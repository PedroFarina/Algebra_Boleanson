<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-62.7917,71.15,33.5083,-37.15</PageViewport>
<gate>
<ID>195</ID>
<type>AA_TOGGLE</type>
<position>-49,13</position>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>196</ID>
<type>AA_TOGGLE</type>
<position>-46,13</position>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_TOGGLE</type>
<position>-41.5,13</position>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_TOGGLE</type>
<position>-38.5,13</position>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>200</ID>
<type>DE_TO</type>
<position>-35.5,32</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>201</ID>
<type>DE_TO</type>
<position>-35.5,29.5</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>202</ID>
<type>DE_TO</type>
<position>-35.5,27</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>203</ID>
<type>DE_TO</type>
<position>-35.5,24.5</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>206</ID>
<type>AA_TOGGLE</type>
<position>-16,13</position>
<output>
<ID>OUT_0</ID>101 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>207</ID>
<type>AA_TOGGLE</type>
<position>-13,13</position>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>211</ID>
<type>DE_TO</type>
<position>-10,27</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>212</ID>
<type>DE_TO</type>
<position>-10,24.5</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>232</ID>
<type>GA_LED</type>
<position>8.5,13</position>
<input>
<ID>N_in3</ID>116 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>233</ID>
<type>GA_LED</type>
<position>12.5,13</position>
<input>
<ID>N_in3</ID>117 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>234</ID>
<type>GA_LED</type>
<position>16.5,13</position>
<input>
<ID>N_in3</ID>118 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>235</ID>
<type>GA_LED</type>
<position>20.5,13</position>
<input>
<ID>N_in3</ID>119 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>239</ID>
<type>DA_FROM</type>
<position>0.5,27</position>
<input>
<ID>IN_0</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID O1</lparam></gate>
<gate>
<ID>240</ID>
<type>DA_FROM</type>
<position>0.5,24.5</position>
<input>
<ID>IN_0</ID>116 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID O0</lparam></gate>
<gate>
<ID>241</ID>
<type>DA_FROM</type>
<position>0.5,29.5</position>
<input>
<ID>IN_0</ID>118 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID O2</lparam></gate>
<gate>
<ID>242</ID>
<type>DA_FROM</type>
<position>0.5,32</position>
<input>
<ID>IN_0</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID O3</lparam></gate>
<gate>
<ID>319</ID>
<type>AA_TOGGLE</type>
<position>-19,13</position>
<output>
<ID>OUT_0</ID>181 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>320</ID>
<type>DE_TO</type>
<position>-10,30</position>
<input>
<ID>IN_0</ID>181 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cin</lparam></gate>
<gate>
<ID>321</ID>
<type>AA_TOGGLE</type>
<position>-22,13</position>
<output>
<ID>OUT_0</ID>182 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>322</ID>
<type>DE_TO</type>
<position>-10,33</position>
<input>
<ID>IN_0</ID>182 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_TOGGLE</type>
<position>-68,13</position>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>162</ID>
<type>AA_TOGGLE</type>
<position>-65,13</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>163</ID>
<type>AA_TOGGLE</type>
<position>-60.5,13</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>164</ID>
<type>AA_TOGGLE</type>
<position>-57.5,13</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>182</ID>
<type>DE_TO</type>
<position>-54.5,32</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>183</ID>
<type>DE_TO</type>
<position>-54.5,29.5</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>184</ID>
<type>DE_TO</type>
<position>-54.5,27</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>185</ID>
<type>DE_TO</type>
<position>-54.5,24.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-57.5,15,-57.5,24.5</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-57.5,24.5,-56.5,24.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>-57.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-60.5,15,-60.5,27</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-60.5,27,-56.5,27</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>-60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-65,15,-65,29.5</points>
<connection>
<GID>162</GID>
<name>OUT_0</name></connection>
<intersection>29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65,29.5,-56.5,29.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>-65 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68,15,-68,32</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68,32,-56.5,32</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>-68 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38.5,15,-38.5,24.5</points>
<connection>
<GID>198</GID>
<name>OUT_0</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-38.5,24.5,-37.5,24.5</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>-38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-41.5,15,-41.5,27</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-41.5,27,-37.5,27</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>-41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,15,-46,29.5</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-46,29.5,-37.5,29.5</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>-46 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,15,-49,32</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<intersection>32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-49,32,-37.5,32</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>-49 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13,15,-13,24.5</points>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,24.5,-12,24.5</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>-13 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,15,-16,27</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,27,-12,27</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,14,8.5,24.5</points>
<connection>
<GID>232</GID>
<name>N_in3</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,24.5,8.5,24.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,14,12.5,27</points>
<connection>
<GID>233</GID>
<name>N_in3</name></connection>
<intersection>27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,27,12.5,27</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,14,16.5,29.5</points>
<connection>
<GID>234</GID>
<name>N_in3</name></connection>
<intersection>29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,29.5,16.5,29.5</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,14,20.5,32</points>
<connection>
<GID>235</GID>
<name>N_in3</name></connection>
<intersection>32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,32,20.5,32</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19,15,-19,30</points>
<connection>
<GID>319</GID>
<name>OUT_0</name></connection>
<intersection>30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-19,30,-12,30</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>-19 0</intersection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,15,-22,33</points>
<connection>
<GID>321</GID>
<name>OUT_0</name></connection>
<intersection>33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-22,33,-12,33</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>-22 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-36.3031,20.2635,116.047,-151.071</PageViewport>
<gate>
<ID>69</ID>
<type>AA_AND2</type>
<position>11,-18.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>AE_OR2</type>
<position>11,-23.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>AI_XOR2</type>
<position>11.5,-33</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>AE_SMALL_INVERTER</type>
<position>10.5,-28.5</position>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_MUX_2x1</type>
<position>31,-22.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>35 </output>
<input>
<ID>SEL_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_MUX_2x1</type>
<position>31,-29.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>36 </output>
<input>
<ID>SEL_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_MUX_2x1</type>
<position>37.5,-26</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>83 </output>
<input>
<ID>SEL_0</ID>82 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>DA_FROM</type>
<position>-16,-10.5</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>90</ID>
<type>DA_FROM</type>
<position>3,-11</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>91</ID>
<type>AA_AND2</type>
<position>11.5,-44.5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>94</ID>
<type>AE_OR2</type>
<position>11.5,-49.5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>AI_XOR2</type>
<position>12,-59</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>96</ID>
<type>AE_SMALL_INVERTER</type>
<position>11,-54.5</position>
<input>
<ID>IN_0</ID>38 </input>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_MUX_2x1</type>
<position>31.5,-48.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>46 </output>
<input>
<ID>SEL_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_MUX_2x1</type>
<position>31.5,-55.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>42 </input>
<output>
<ID>OUT</ID>47 </output>
<input>
<ID>SEL_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_MUX_2x1</type>
<position>38,-52</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>84 </output>
<input>
<ID>SEL_0</ID>82 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>101</ID>
<type>DA_FROM</type>
<position>-19.5,-10.5</position>
<input>
<ID>IN_0</ID>38 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>102</ID>
<type>DA_FROM</type>
<position>-0.5,-11</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_AND2</type>
<position>12.5,-70.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AE_OR2</type>
<position>12.5,-75.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>AI_XOR2</type>
<position>13,-85</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>AE_SMALL_INVERTER</type>
<position>12,-80.5</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_MUX_2x1</type>
<position>32.5,-74.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>57 </output>
<input>
<ID>SEL_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_MUX_2x1</type>
<position>32.5,-81.5</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>58 </output>
<input>
<ID>SEL_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_MUX_2x1</type>
<position>39,-78</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>85 </output>
<input>
<ID>SEL_0</ID>82 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>DA_FROM</type>
<position>-23.5,-10.5</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>114</ID>
<type>DA_FROM</type>
<position>-4.5,-11</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_AND2</type>
<position>13,-97</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AE_OR2</type>
<position>13,-102</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>AI_XOR2</type>
<position>13.5,-111.5</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AE_SMALL_INVERTER</type>
<position>12.5,-107</position>
<input>
<ID>IN_0</ID>60 </input>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_MUX_2x1</type>
<position>33,-101</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>68 </output>
<input>
<ID>SEL_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_MUX_2x1</type>
<position>33,-108</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>69 </output>
<input>
<ID>SEL_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_MUX_2x1</type>
<position>39.5,-104.5</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>86 </output>
<input>
<ID>SEL_0</ID>82 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>-27,-10.5</position>
<input>
<ID>IN_0</ID>60 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>126</ID>
<type>DA_FROM</type>
<position>-8,-11</position>
<input>
<ID>IN_0</ID>61 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>139</ID>
<type>DA_FROM</type>
<position>26.5,-10.5</position>
<input>
<ID>IN_0</ID>40 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>140</ID>
<type>DA_FROM</type>
<position>34,-10.5</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>142</ID>
<type>DE_TO</type>
<position>44.5,-10.5</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O3</lparam></gate>
<gate>
<ID>143</ID>
<type>DE_TO</type>
<position>48.5,-10.5</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O2</lparam></gate>
<gate>
<ID>144</ID>
<type>DE_TO</type>
<position>52,-10.5</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O1</lparam></gate>
<gate>
<ID>145</ID>
<type>DE_TO</type>
<position>55,-10.5</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID O0</lparam></gate>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-34,-16,-12.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>-34 3</intersection>
<intersection>-28.5 8</intersection>
<intersection>-24.5 5</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-19.5,8,-19.5</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-16,-34,8.5,-34</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-16,-24.5,8,-24.5</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-16,-28.5,8.5,-28.5</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-32,3,-13</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>-32 3</intersection>
<intersection>-22.5 4</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,-17.5,8,-17.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>3,-32,8.5,-32</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>3,-22.5,8,-22.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-33,21.5,-30.5</points>
<intersection>-33 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-30.5,29,-30.5</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-33,21.5,-33</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,-28.5,29,-28.5</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<connection>
<GID>84</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14,-23.5,29,-23.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<connection>
<GID>77</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-21.5,21.5,-18.5</points>
<intersection>-21.5 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-21.5,29,-21.5</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-18.5,21.5,-18.5</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-25,34,-22.5</points>
<intersection>-25 1</intersection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-25,35.5,-25</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-22.5,34,-22.5</points>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-29.5,34,-27</points>
<intersection>-29.5 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-27,35.5,-27</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-29.5,34,-29.5</points>
<connection>
<GID>84</GID>
<name>OUT</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,-60,-19.5,-12.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-60 3</intersection>
<intersection>-54.5 8</intersection>
<intersection>-50.5 5</intersection>
<intersection>-45.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-19.5,-45.5,8.5,-45.5</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-19.5,-60,9,-60</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-19.5,-50.5,8.5,-50.5</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-19.5,-54.5,9,-54.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>-19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,-58,-0.5,-13</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>-58 3</intersection>
<intersection>-48.5 4</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-0.5,-43.5,8.5,-43.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>-0.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-0.5,-58,9,-58</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>-0.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-0.5,-48.5,8.5,-48.5</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>-0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-105.5,26.5,-12.5</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>-105.5 28</intersection>
<intersection>-97.5 29</intersection>
<intersection>-79 20</intersection>
<intersection>-71 21</intersection>
<intersection>-53 4</intersection>
<intersection>-45 5</intersection>
<intersection>-27 12</intersection>
<intersection>-19 13</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>26.5,-53,31.5,-53</points>
<connection>
<GID>98</GID>
<name>SEL_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>26.5,-45,31.5,-45</points>
<intersection>26.5 0</intersection>
<intersection>31.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>31.5,-46,31.5,-45</points>
<connection>
<GID>97</GID>
<name>SEL_0</name></connection>
<intersection>-45 5</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>26.5,-27,31,-27</points>
<connection>
<GID>84</GID>
<name>SEL_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>26.5,-19,31,-19</points>
<intersection>26.5 0</intersection>
<intersection>31 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>31,-20,31,-19</points>
<connection>
<GID>83</GID>
<name>SEL_0</name></connection>
<intersection>-19 13</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>26.5,-79,32.5,-79</points>
<connection>
<GID>110</GID>
<name>SEL_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>26.5,-71,32.5,-71</points>
<intersection>26.5 0</intersection>
<intersection>32.5 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>32.5,-72,32.5,-71</points>
<connection>
<GID>109</GID>
<name>SEL_0</name></connection>
<intersection>-71 21</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>26.5,-105.5,33,-105.5</points>
<connection>
<GID>122</GID>
<name>SEL_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>26.5,-97.5,33,-97.5</points>
<intersection>26.5 0</intersection>
<intersection>33 30</intersection></hsegment>
<vsegment>
<ID>30</ID>
<points>33,-98.5,33,-97.5</points>
<connection>
<GID>121</GID>
<name>SEL_0</name></connection>
<intersection>-97.5 29</intersection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-59,22,-56.5</points>
<intersection>-59 2</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-56.5,29.5,-56.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,-59,22,-59</points>
<connection>
<GID>95</GID>
<name>OUT</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-54.5,29.5,-54.5</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14.5,-49.5,29.5,-49.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<connection>
<GID>94</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22,-47.5,22,-44.5</points>
<intersection>-47.5 1</intersection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-47.5,29.5,-47.5</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<intersection>22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-44.5,22,-44.5</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<intersection>22 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-51,34.5,-48.5</points>
<intersection>-51 1</intersection>
<intersection>-48.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-51,36,-51</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,-48.5,34.5,-48.5</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-55.5,34.5,-53</points>
<intersection>-55.5 2</intersection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-53,36,-53</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,-55.5,34.5,-55.5</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-23.5,-86,-23.5,-12.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>-86 3</intersection>
<intersection>-80.5 8</intersection>
<intersection>-76.5 5</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-23.5,-71.5,9.5,-71.5</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>-23.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-23.5,-86,10,-86</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>-23.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-23.5,-76.5,9.5,-76.5</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>-23.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-23.5,-80.5,10,-80.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-84,-4.5,-13</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>-84 3</intersection>
<intersection>-74.5 4</intersection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-69.5,9.5,-69.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-4.5,-84,10,-84</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-4.5,-74.5,9.5,-74.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-85,23,-82.5</points>
<intersection>-85 2</intersection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-82.5,30.5,-82.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-85,23,-85</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14,-80.5,30.5,-80.5</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<connection>
<GID>110</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15.5,-75.5,30.5,-75.5</points>
<connection>
<GID>106</GID>
<name>OUT</name></connection>
<connection>
<GID>109</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-73.5,23,-70.5</points>
<intersection>-73.5 1</intersection>
<intersection>-70.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-73.5,30.5,-73.5</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15.5,-70.5,23,-70.5</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-77,35.5,-74.5</points>
<intersection>-77 1</intersection>
<intersection>-74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-77,37,-77</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-74.5,35.5,-74.5</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-81.5,35.5,-79</points>
<intersection>-81.5 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-79,37,-79</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-81.5,35.5,-81.5</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27,-112.5,-27,-12.5</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>-112.5 3</intersection>
<intersection>-107 8</intersection>
<intersection>-103 5</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27,-98,10,-98</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<intersection>-27 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-27,-112.5,10.5,-112.5</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>-27 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-27,-103,10,-103</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>-27 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-27,-107,10.5,-107</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>-27 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,-110.5,-8,-13</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>-110.5 3</intersection>
<intersection>-101 4</intersection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8,-96,10,-96</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>-8 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-8,-110.5,10.5,-110.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-8 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-8,-101,10,-101</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>-8 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-111.5,23.5,-109</points>
<intersection>-111.5 2</intersection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-109,31,-109</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-111.5,23.5,-111.5</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14.5,-107,31,-107</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-102,31,-102</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<connection>
<GID>118</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-100,23.5,-97</points>
<intersection>-100 1</intersection>
<intersection>-97 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-100,31,-100</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-97,23.5,-97</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-103.5,36,-101</points>
<intersection>-103.5 1</intersection>
<intersection>-101 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-103.5,37.5,-103.5</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-101,36,-101</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-108,36,-105.5</points>
<intersection>-108 2</intersection>
<intersection>-105.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-105.5,37.5,-105.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-108,36,-108</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-97.5,34,-12.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>-97.5 5</intersection>
<intersection>-73 6</intersection>
<intersection>-47 3</intersection>
<intersection>-21 7</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>34,-47,38,-47</points>
<intersection>34 0</intersection>
<intersection>38 8</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>34,-97.5,39.5,-97.5</points>
<intersection>34 0</intersection>
<intersection>39.5 11</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>34,-73,39,-73</points>
<intersection>34 0</intersection>
<intersection>39 10</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>34,-21,37.5,-21</points>
<intersection>34 0</intersection>
<intersection>37.5 9</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>38,-49.5,38,-47</points>
<connection>
<GID>99</GID>
<name>SEL_0</name></connection>
<intersection>-47 3</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>37.5,-23.5,37.5,-21</points>
<connection>
<GID>85</GID>
<name>SEL_0</name></connection>
<intersection>-21 7</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>39,-75.5,39,-73</points>
<connection>
<GID>111</GID>
<name>SEL_0</name></connection>
<intersection>-73 6</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>39.5,-102,39.5,-97.5</points>
<connection>
<GID>123</GID>
<name>SEL_0</name></connection>
<intersection>-97.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-26,55,-12.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-26,55,-26</points>
<connection>
<GID>85</GID>
<name>OUT</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-52,52,-12.5</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>-52 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-52,52,-52</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48.5,-78,48.5,-12.5</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-78,48.5,-78</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<intersection>48.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-104.5,44.5,-12.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>-104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-104.5,44.5,-104.5</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-36.6403,14.5271,59.6597,-93.7729</PageViewport>
<gate>
<ID>601</ID>
<type>DA_FROM</type>
<position>48,-17.5</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Si0</lparam></gate>
<gate>
<ID>602</ID>
<type>DA_FROM</type>
<position>48.5,-31</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Si0</lparam></gate>
<gate>
<ID>603</ID>
<type>DA_FROM</type>
<position>48,-44</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Si0</lparam></gate>
<gate>
<ID>604</ID>
<type>DA_FROM</type>
<position>48,-59</position>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Si0</lparam></gate>
<gate>
<ID>243</ID>
<type>DA_FROM</type>
<position>-17.5,-5.5</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>244</ID>
<type>DA_FROM</type>
<position>1.5,-6</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B0</lparam></gate>
<gate>
<ID>245</ID>
<type>DA_FROM</type>
<position>-21,-5.5</position>
<input>
<ID>IN_0</ID>128 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>246</ID>
<type>DA_FROM</type>
<position>-2,-6</position>
<input>
<ID>IN_0</ID>126 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>247</ID>
<type>DA_FROM</type>
<position>-25,-5.5</position>
<input>
<ID>IN_0</ID>132 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>248</ID>
<type>DA_FROM</type>
<position>-6,-6</position>
<input>
<ID>IN_0</ID>130 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>249</ID>
<type>DA_FROM</type>
<position>-28.5,-5.5</position>
<input>
<ID>IN_0</ID>136 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>250</ID>
<type>DA_FROM</type>
<position>-9.5,-6</position>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_MUX_2x1</type>
<position>25.5,-14</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>122 </input>
<output>
<ID>OUT</ID>144 </output>
<input>
<ID>SEL_0</ID>121 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_MUX_2x1</type>
<position>25.5,-20.5</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>122 </input>
<output>
<ID>OUT</ID>143 </output>
<input>
<ID>SEL_0</ID>121 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>256</ID>
<type>DA_FROM</type>
<position>9,-5.5</position>
<input>
<ID>IN_0</ID>121 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>257</ID>
<type>DA_FROM</type>
<position>29,-7</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>259</ID>
<type>AE_SMALL_INVERTER</type>
<position>20.5,-15</position>
<input>
<ID>IN_0</ID>124 </input>
<output>
<ID>OUT_0</ID>123 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>260</ID>
<type>AA_MUX_2x1</type>
<position>25.5,-28</position>
<input>
<ID>IN_0</ID>127 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>142 </output>
<input>
<ID>SEL_0</ID>121 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>261</ID>
<type>AA_MUX_2x1</type>
<position>25.5,-34.5</position>
<input>
<ID>IN_0</ID>128 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>141 </output>
<input>
<ID>SEL_0</ID>121 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>262</ID>
<type>AE_SMALL_INVERTER</type>
<position>20.5,-29</position>
<input>
<ID>IN_0</ID>128 </input>
<output>
<ID>OUT_0</ID>127 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>263</ID>
<type>AA_MUX_2x1</type>
<position>25,-41.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>140 </output>
<input>
<ID>SEL_0</ID>121 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_MUX_2x1</type>
<position>25,-48</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>139 </output>
<input>
<ID>SEL_0</ID>121 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>265</ID>
<type>AE_SMALL_INVERTER</type>
<position>20,-42.5</position>
<input>
<ID>IN_0</ID>132 </input>
<output>
<ID>OUT_0</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>266</ID>
<type>AA_MUX_2x1</type>
<position>25,-56</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>134 </input>
<output>
<ID>OUT</ID>138 </output>
<input>
<ID>SEL_0</ID>121 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>267</ID>
<type>AA_MUX_2x1</type>
<position>25,-62.5</position>
<input>
<ID>IN_0</ID>136 </input>
<input>
<ID>IN_1</ID>134 </input>
<output>
<ID>OUT</ID>137 </output>
<input>
<ID>SEL_0</ID>121 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>268</ID>
<type>AE_SMALL_INVERTER</type>
<position>20,-57</position>
<input>
<ID>IN_0</ID>136 </input>
<output>
<ID>OUT_0</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>269</ID>
<type>AA_MUX_2x1</type>
<position>31.5,-17.5</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>144 </input>
<output>
<ID>OUT</ID>146 </output>
<input>
<ID>SEL_0</ID>145 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>270</ID>
<type>AA_MUX_2x1</type>
<position>31.5,-31</position>
<input>
<ID>IN_0</ID>141 </input>
<input>
<ID>IN_1</ID>142 </input>
<output>
<ID>OUT</ID>147 </output>
<input>
<ID>SEL_0</ID>145 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>271</ID>
<type>AA_MUX_2x1</type>
<position>31,-44.5</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>140 </input>
<output>
<ID>OUT</ID>148 </output>
<input>
<ID>SEL_0</ID>145 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>272</ID>
<type>AA_MUX_2x1</type>
<position>31.5,-59</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>149 </output>
<input>
<ID>SEL_0</ID>145 </input>
<gparam>angle 0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>276</ID>
<type>DE_TO</type>
<position>37,-17.5</position>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M0</lparam></gate>
<gate>
<ID>277</ID>
<type>DE_TO</type>
<position>36.5,-31</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M1</lparam></gate>
<gate>
<ID>278</ID>
<type>DE_TO</type>
<position>36,-44.5</position>
<input>
<ID>IN_0</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M2</lparam></gate>
<gate>
<ID>279</ID>
<type>DE_TO</type>
<position>36.5,-59</position>
<input>
<ID>IN_0</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M3</lparam></gate>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-32,9,-7.5</points>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>-32 12</intersection>
<intersection>-24 13</intersection>
<intersection>-18 4</intersection>
<intersection>-10 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>9,-18,25.5,-18</points>
<connection>
<GID>255</GID>
<name>SEL_0</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>9,-10,25.5,-10</points>
<intersection>9 0</intersection>
<intersection>25.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>25.5,-11.5,25.5,-10</points>
<connection>
<GID>254</GID>
<name>SEL_0</name></connection>
<intersection>-10 5</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>8.5,-32,25.5,-32</points>
<connection>
<GID>261</GID>
<name>SEL_0</name></connection>
<intersection>8.5 15</intersection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>9,-24,25.5,-24</points>
<intersection>9 0</intersection>
<intersection>25.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>25.5,-25.5,25.5,-24</points>
<connection>
<GID>260</GID>
<name>SEL_0</name></connection>
<intersection>-24 13</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>8.5,-60,8.5,-32</points>
<intersection>-60 28</intersection>
<intersection>-52 29</intersection>
<intersection>-45.5 20</intersection>
<intersection>-37.5 21</intersection>
<intersection>-32 12</intersection></vsegment>
<hsegment>
<ID>20</ID>
<points>8.5,-45.5,25,-45.5</points>
<connection>
<GID>264</GID>
<name>SEL_0</name></connection>
<intersection>8.5 15</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>8.5,-37.5,25,-37.5</points>
<intersection>8.5 15</intersection>
<intersection>25 22</intersection></hsegment>
<vsegment>
<ID>22</ID>
<points>25,-39,25,-37.5</points>
<connection>
<GID>263</GID>
<name>SEL_0</name></connection>
<intersection>-37.5 21</intersection></vsegment>
<hsegment>
<ID>28</ID>
<points>8.5,-60,25,-60</points>
<connection>
<GID>267</GID>
<name>SEL_0</name></connection>
<intersection>8.5 15</intersection></hsegment>
<hsegment>
<ID>29</ID>
<points>8.5,-52,25,-52</points>
<intersection>8.5 15</intersection>
<intersection>25 30</intersection></hsegment>
<vsegment>
<ID>30</ID>
<points>25,-53.5,25,-52</points>
<connection>
<GID>266</GID>
<name>SEL_0</name></connection>
<intersection>-52 29</intersection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1.5,-19.5,1.5,-8</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>-19.5 3</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1.5,-13,23.5,-13</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<intersection>1.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>1.5,-19.5,23.5,-19.5</points>
<connection>
<GID>255</GID>
<name>IN_1</name></connection>
<intersection>1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-15,23.5,-15</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<connection>
<GID>259</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-17.5,-21.5,-17.5,-7.5</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>-21.5 3</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-17.5,-15,18.5,-15</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<intersection>-17.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-17.5,-21.5,23.5,-21.5</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>-17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2,-33.5,-2,-8</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>-33.5 3</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2,-27,23.5,-27</points>
<connection>
<GID>260</GID>
<name>IN_1</name></connection>
<intersection>-2 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-2,-33.5,23.5,-33.5</points>
<connection>
<GID>261</GID>
<name>IN_1</name></connection>
<intersection>-2 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22.5,-29,23.5,-29</points>
<connection>
<GID>262</GID>
<name>OUT_0</name></connection>
<connection>
<GID>260</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-21,-35.5,-21,-7.5</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>-35.5 3</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-21,-29,18.5,-29</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>-21 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-21,-35.5,23.5,-35.5</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>-21 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6,-47,-6,-8</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>-47 3</intersection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6,-40.5,23,-40.5</points>
<connection>
<GID>263</GID>
<name>IN_1</name></connection>
<intersection>-6 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-6,-47,23,-47</points>
<connection>
<GID>264</GID>
<name>IN_1</name></connection>
<intersection>-6 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-42.5,23,-42.5</points>
<connection>
<GID>265</GID>
<name>OUT_0</name></connection>
<connection>
<GID>263</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25,-49,-25,-7.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>-49 3</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25,-42.5,18,-42.5</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>-25 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-25,-49,23,-49</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>-25 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-9.5,-61.5,-9.5,-8</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>-61.5 3</intersection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-9.5,-55,23,-55</points>
<connection>
<GID>266</GID>
<name>IN_1</name></connection>
<intersection>-9.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-9.5,-61.5,23,-61.5</points>
<connection>
<GID>267</GID>
<name>IN_1</name></connection>
<intersection>-9.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-57,23,-57</points>
<connection>
<GID>268</GID>
<name>OUT_0</name></connection>
<connection>
<GID>266</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28.5,-63.5,-28.5,-7.5</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>-63.5 3</intersection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-28.5,-57,18,-57</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>-28.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-28.5,-63.5,23,-63.5</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>-28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-62.5,28,-60</points>
<intersection>-62.5 1</intersection>
<intersection>-60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-62.5,28,-62.5</points>
<connection>
<GID>267</GID>
<name>OUT</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-60,29.5,-60</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-58,28,-56</points>
<intersection>-58 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-56,28,-56</points>
<connection>
<GID>266</GID>
<name>OUT</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-58,29.5,-58</points>
<connection>
<GID>272</GID>
<name>IN_1</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-48,28,-45.5</points>
<intersection>-48 1</intersection>
<intersection>-45.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-48,28,-48</points>
<connection>
<GID>264</GID>
<name>OUT</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-45.5,29,-45.5</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-43.5,28,-41.5</points>
<intersection>-43.5 2</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-41.5,28,-41.5</points>
<connection>
<GID>263</GID>
<name>OUT</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-43.5,29,-43.5</points>
<connection>
<GID>271</GID>
<name>IN_1</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-34.5,28.5,-32</points>
<intersection>-34.5 1</intersection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-34.5,28.5,-34.5</points>
<connection>
<GID>261</GID>
<name>OUT</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-32,29.5,-32</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-30,28.5,-28</points>
<intersection>-30 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-28,28.5,-28</points>
<connection>
<GID>260</GID>
<name>OUT</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-30,29.5,-30</points>
<connection>
<GID>270</GID>
<name>IN_1</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-20.5,28.5,-18.5</points>
<intersection>-20.5 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-20.5,28.5,-20.5</points>
<connection>
<GID>255</GID>
<name>OUT</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-18.5,29.5,-18.5</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-16.5,28.5,-14</points>
<intersection>-16.5 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-14,28.5,-14</points>
<connection>
<GID>254</GID>
<name>OUT</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-16.5,29.5,-16.5</points>
<connection>
<GID>269</GID>
<name>IN_1</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-56.5,29,-9</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>-56.5 6</intersection>
<intersection>-42 4</intersection>
<intersection>-28.5 7</intersection>
<intersection>-15 8</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>29,-42,31,-42</points>
<connection>
<GID>271</GID>
<name>SEL_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>29,-56.5,31.5,-56.5</points>
<connection>
<GID>272</GID>
<name>SEL_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>29,-28.5,31.5,-28.5</points>
<connection>
<GID>270</GID>
<name>SEL_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>29,-15,31.5,-15</points>
<connection>
<GID>269</GID>
<name>SEL_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-17.5,35,-17.5</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>33.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33.5,-17.5,33.5,-17.5</points>
<connection>
<GID>269</GID>
<name>OUT</name></connection>
<intersection>-17.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-31,34.5,-31</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>33.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33.5,-31,33.5,-31</points>
<connection>
<GID>270</GID>
<name>OUT</name></connection>
<intersection>-31 1</intersection></vsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33,-44.5,34,-44.5</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>33 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33,-44.5,33,-44.5</points>
<connection>
<GID>271</GID>
<name>OUT</name></connection>
<intersection>-44.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-59,34.5,-59</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<intersection>33.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33.5,-59,33.5,-59</points>
<connection>
<GID>272</GID>
<name>OUT</name></connection>
<intersection>-59 1</intersection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>-542.696,108.445,-457,12.0692</PageViewport>
<gate>
<ID>386</ID>
<type>DA_FROM</type>
<position>-565,104.5</position>
<input>
<ID>IN_0</ID>207 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M1</lparam></gate>
<gate>
<ID>387</ID>
<type>DA_FROM</type>
<position>-566,76.5</position>
<input>
<ID>IN_0</ID>221 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>388</ID>
<type>DA_FROM</type>
<position>-565,71.5</position>
<input>
<ID>IN_0</ID>220 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M2</lparam></gate>
<gate>
<ID>389</ID>
<type>DA_FROM</type>
<position>-565.5,44.5</position>
<input>
<ID>IN_0</ID>234 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>390</ID>
<type>DA_FROM</type>
<position>-564.5,39</position>
<input>
<ID>IN_0</ID>233 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M3</lparam></gate>
<gate>
<ID>281</ID>
<type>BA_NAND2</type>
<position>-553.5,137.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>156 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>282</ID>
<type>BA_NAND2</type>
<position>-539.5,141</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>158 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>283</ID>
<type>BA_NAND2</type>
<position>-539.5,134</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>156 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>284</ID>
<type>BA_NAND2</type>
<position>-527.5,137</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>154 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>285</ID>
<type>BA_NAND2</type>
<position>-514,141</position>
<input>
<ID>IN_0</ID>152 </input>
<input>
<ID>IN_1</ID>153 </input>
<output>
<ID>OUT</ID>150 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>286</ID>
<type>BA_NAND2</type>
<position>-502.5,145</position>
<input>
<ID>IN_0</ID>152 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>287</ID>
<type>BA_NAND2</type>
<position>-502.5,137</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>153 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>288</ID>
<type>BA_NAND2</type>
<position>-490.5,141</position>
<input>
<ID>IN_0</ID>160 </input>
<input>
<ID>IN_1</ID>159 </input>
<output>
<ID>OUT</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>289</ID>
<type>BA_NAND2</type>
<position>-502.5,124.5</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>158 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>293</ID>
<type>DA_FROM</type>
<position>-564.5,140</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>294</ID>
<type>DA_FROM</type>
<position>-563.5,135</position>
<input>
<ID>IN_0</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M0</lparam></gate>
<gate>
<ID>317</ID>
<type>DA_FROM</type>
<position>-571,160.5</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>318</ID>
<type>DA_FROM</type>
<position>-567.5,160.5</position>
<input>
<ID>IN_0</ID>184 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>323</ID>
<type>DA_FROM</type>
<position>-556,160.5</position>
<input>
<ID>IN_0</ID>186 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Cin</lparam></gate>
<gate>
<ID>325</ID>
<type>AI_XOR2</type>
<position>-561.5,149.5</position>
<input>
<ID>IN_0</ID>184 </input>
<input>
<ID>IN_1</ID>183 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>327</ID>
<type>AA_AND2</type>
<position>-549.5,150.5</position>
<input>
<ID>IN_0</ID>186 </input>
<input>
<ID>IN_1</ID>185 </input>
<output>
<ID>OUT</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>329</ID>
<type>DE_TO</type>
<position>-483,141</position>
<input>
<ID>IN_0</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Si0</lparam></gate>
<gate>
<ID>330</ID>
<type>DE_TO</type>
<position>-494.5,124.5</position>
<input>
<ID>IN_0</ID>203 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cout0</lparam></gate>
<gate>
<ID>344</ID>
<type>BA_NAND2</type>
<position>-553.5,107</position>
<input>
<ID>IN_0</ID>208 </input>
<input>
<ID>IN_1</ID>207 </input>
<output>
<ID>OUT</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>345</ID>
<type>BA_NAND2</type>
<position>-539.5,110.5</position>
<input>
<ID>IN_0</ID>208 </input>
<input>
<ID>IN_1</ID>209 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>346</ID>
<type>BA_NAND2</type>
<position>-539.5,103.5</position>
<input>
<ID>IN_0</ID>209 </input>
<input>
<ID>IN_1</ID>207 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>347</ID>
<type>BA_NAND2</type>
<position>-527.5,106.5</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>205 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>348</ID>
<type>BA_NAND2</type>
<position>-514,110.5</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>204 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>349</ID>
<type>BA_NAND2</type>
<position>-502.5,114.5</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>202 </input>
<output>
<ID>OUT</ID>211 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>350</ID>
<type>BA_NAND2</type>
<position>-502.5,106.5</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>204 </input>
<output>
<ID>OUT</ID>210 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>351</ID>
<type>BA_NAND2</type>
<position>-490.5,110.5</position>
<input>
<ID>IN_0</ID>211 </input>
<input>
<ID>IN_1</ID>210 </input>
<output>
<ID>OUT</ID>213 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>352</ID>
<type>BA_NAND2</type>
<position>-502.5,94</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>209 </input>
<output>
<ID>OUT</ID>216 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>355</ID>
<type>DE_TO</type>
<position>-483,110.5</position>
<input>
<ID>IN_0</ID>213 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Si1</lparam></gate>
<gate>
<ID>356</ID>
<type>DE_TO</type>
<position>-494.5,94</position>
<input>
<ID>IN_0</ID>216 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cout1</lparam></gate>
<gate>
<ID>357</ID>
<type>BA_NAND2</type>
<position>-553,74.5</position>
<input>
<ID>IN_0</ID>221 </input>
<input>
<ID>IN_1</ID>220 </input>
<output>
<ID>OUT</ID>222 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>358</ID>
<type>BA_NAND2</type>
<position>-539,78</position>
<input>
<ID>IN_0</ID>221 </input>
<input>
<ID>IN_1</ID>222 </input>
<output>
<ID>OUT</ID>219 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>359</ID>
<type>BA_NAND2</type>
<position>-539,71</position>
<input>
<ID>IN_0</ID>222 </input>
<input>
<ID>IN_1</ID>220 </input>
<output>
<ID>OUT</ID>218 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>360</ID>
<type>BA_NAND2</type>
<position>-527,74</position>
<input>
<ID>IN_0</ID>219 </input>
<input>
<ID>IN_1</ID>218 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>BA_NAND2</type>
<position>-513.5,78</position>
<input>
<ID>IN_0</ID>216 </input>
<input>
<ID>IN_1</ID>217 </input>
<output>
<ID>OUT</ID>215 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>362</ID>
<type>BA_NAND2</type>
<position>-502,82</position>
<input>
<ID>IN_0</ID>216 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>363</ID>
<type>BA_NAND2</type>
<position>-502,74</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>217 </input>
<output>
<ID>OUT</ID>223 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>364</ID>
<type>BA_NAND2</type>
<position>-490,78</position>
<input>
<ID>IN_0</ID>224 </input>
<input>
<ID>IN_1</ID>223 </input>
<output>
<ID>OUT</ID>226 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>365</ID>
<type>BA_NAND2</type>
<position>-502,61.5</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>222 </input>
<output>
<ID>OUT</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>368</ID>
<type>DE_TO</type>
<position>-482.5,78</position>
<input>
<ID>IN_0</ID>226 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Si2</lparam></gate>
<gate>
<ID>369</ID>
<type>DE_TO</type>
<position>-494,61.5</position>
<input>
<ID>IN_0</ID>229 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cout2</lparam></gate>
<gate>
<ID>370</ID>
<type>BA_NAND2</type>
<position>-553,41.5</position>
<input>
<ID>IN_0</ID>234 </input>
<input>
<ID>IN_1</ID>233 </input>
<output>
<ID>OUT</ID>235 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>371</ID>
<type>BA_NAND2</type>
<position>-539,45</position>
<input>
<ID>IN_0</ID>234 </input>
<input>
<ID>IN_1</ID>235 </input>
<output>
<ID>OUT</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>372</ID>
<type>BA_NAND2</type>
<position>-539,38</position>
<input>
<ID>IN_0</ID>235 </input>
<input>
<ID>IN_1</ID>233 </input>
<output>
<ID>OUT</ID>231 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>373</ID>
<type>BA_NAND2</type>
<position>-527,41</position>
<input>
<ID>IN_0</ID>232 </input>
<input>
<ID>IN_1</ID>231 </input>
<output>
<ID>OUT</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>374</ID>
<type>BA_NAND2</type>
<position>-513.5,45</position>
<input>
<ID>IN_0</ID>229 </input>
<input>
<ID>IN_1</ID>230 </input>
<output>
<ID>OUT</ID>228 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>375</ID>
<type>BA_NAND2</type>
<position>-502,49</position>
<input>
<ID>IN_0</ID>229 </input>
<input>
<ID>IN_1</ID>228 </input>
<output>
<ID>OUT</ID>237 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>376</ID>
<type>BA_NAND2</type>
<position>-502,41</position>
<input>
<ID>IN_0</ID>228 </input>
<input>
<ID>IN_1</ID>230 </input>
<output>
<ID>OUT</ID>236 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>377</ID>
<type>BA_NAND2</type>
<position>-490,45</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>236 </input>
<output>
<ID>OUT</ID>239 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>378</ID>
<type>BA_NAND2</type>
<position>-502,28.5</position>
<input>
<ID>IN_0</ID>228 </input>
<input>
<ID>IN_1</ID>235 </input>
<output>
<ID>OUT</ID>240 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>381</ID>
<type>DE_TO</type>
<position>-482.5,45</position>
<input>
<ID>IN_0</ID>239 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Si3</lparam></gate>
<gate>
<ID>382</ID>
<type>DE_TO</type>
<position>-494,28.5</position>
<input>
<ID>IN_0</ID>240 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cout3</lparam></gate>
<gate>
<ID>385</ID>
<type>DA_FROM</type>
<position>-566,109.5</position>
<input>
<ID>IN_0</ID>208 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-506.5,95,-506.5,113.5</points>
<intersection>95 2</intersection>
<intersection>110.5 3</intersection>
<intersection>113.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-506.5,113.5,-505.5,113.5</points>
<connection>
<GID>349</GID>
<name>IN_1</name></connection>
<intersection>-506.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-506.5,95,-505.5,95</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>-506.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-511,110.5,-506.5,110.5</points>
<connection>
<GID>348</GID>
<name>OUT</name></connection>
<intersection>-508 4</intersection>
<intersection>-506.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-508,107.5,-508,110.5</points>
<intersection>107.5 6</intersection>
<intersection>110.5 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-508,107.5,-505.5,107.5</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<intersection>-508 4</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-519,111.5,-519,115.5</points>
<intersection>111.5 2</intersection>
<intersection>115.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-519,115.5,-505.5,115.5</points>
<connection>
<GID>349</GID>
<name>IN_0</name></connection>
<intersection>-519 0</intersection>
<intersection>-509 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-519,111.5,-517,111.5</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<intersection>-519 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-509,115.5,-509,124.5</points>
<intersection>115.5 1</intersection>
<intersection>124.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-509,124.5,-496.5,124.5</points>
<connection>
<GID>289</GID>
<name>OUT</name></connection>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>-509 3</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-519,105.5,-519,109.5</points>
<intersection>105.5 2</intersection>
<intersection>106.5 3</intersection>
<intersection>109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-519,109.5,-517,109.5</points>
<connection>
<GID>348</GID>
<name>IN_1</name></connection>
<intersection>-519 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-519,105.5,-505.5,105.5</points>
<connection>
<GID>350</GID>
<name>IN_1</name></connection>
<intersection>-519 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-524.5,106.5,-519,106.5</points>
<connection>
<GID>347</GID>
<name>OUT</name></connection>
<intersection>-519 0</intersection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-533.5,103.5,-533.5,105.5</points>
<intersection>103.5 2</intersection>
<intersection>105.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-533.5,105.5,-530.5,105.5</points>
<connection>
<GID>347</GID>
<name>IN_1</name></connection>
<intersection>-533.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-536.5,103.5,-533.5,103.5</points>
<connection>
<GID>346</GID>
<name>OUT</name></connection>
<intersection>-533.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-533.5,107.5,-533.5,110.5</points>
<intersection>107.5 1</intersection>
<intersection>110.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-533.5,107.5,-530.5,107.5</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>-533.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-536.5,110.5,-533.5,110.5</points>
<connection>
<GID>345</GID>
<name>OUT</name></connection>
<intersection>-533.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-559,102.5,-542.5,102.5</points>
<connection>
<GID>346</GID>
<name>IN_1</name></connection>
<intersection>-559 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-559,102.5,-559,104.5</points>
<intersection>102.5 1</intersection>
<intersection>104.5 6</intersection>
<intersection>104.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-563,104.5,-556.5,104.5</points>
<connection>
<GID>386</GID>
<name>IN_0</name></connection>
<intersection>-559 4</intersection>
<intersection>-556.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-556.5,104.5,-556.5,106</points>
<connection>
<GID>344</GID>
<name>IN_1</name></connection>
<intersection>104.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-559,111.5,-542.5,111.5</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<intersection>-559 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-559,109.5,-559,111.5</points>
<intersection>109.5 6</intersection>
<intersection>109.5 6</intersection>
<intersection>111.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-564,109.5,-556.5,109.5</points>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>-559 4</intersection>
<intersection>-556.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-556.5,108,-556.5,109.5</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>109.5 6</intersection></vsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-546.5,93,-546.5,109.5</points>
<intersection>93 3</intersection>
<intersection>104.5 6</intersection>
<intersection>107 1</intersection>
<intersection>109.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-550.5,107,-546.5,107</points>
<connection>
<GID>344</GID>
<name>OUT</name></connection>
<intersection>-546.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-546.5,109.5,-542.5,109.5</points>
<connection>
<GID>345</GID>
<name>IN_1</name></connection>
<intersection>-546.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-546.5,93,-505.5,93</points>
<connection>
<GID>352</GID>
<name>IN_1</name></connection>
<intersection>-546.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-546.5,104.5,-542.5,104.5</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>-546.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-496.5,106.5,-496.5,109.5</points>
<intersection>106.5 2</intersection>
<intersection>109.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-496.5,109.5,-493.5,109.5</points>
<connection>
<GID>351</GID>
<name>IN_1</name></connection>
<intersection>-496.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-499.5,106.5,-496.5,106.5</points>
<connection>
<GID>350</GID>
<name>OUT</name></connection>
<intersection>-496.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-496.5,111.5,-496.5,114.5</points>
<intersection>111.5 1</intersection>
<intersection>114.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-496.5,111.5,-493.5,111.5</points>
<connection>
<GID>351</GID>
<name>IN_0</name></connection>
<intersection>-496.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-499.5,114.5,-496.5,114.5</points>
<connection>
<GID>349</GID>
<name>OUT</name></connection>
<intersection>-496.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-487.5,110.5,-485,110.5</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>-487.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-487.5,110.5,-487.5,110.5</points>
<connection>
<GID>351</GID>
<name>OUT</name></connection>
<intersection>110.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-506,62.5,-506,81</points>
<intersection>62.5 2</intersection>
<intersection>78 3</intersection>
<intersection>81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-506,81,-505,81</points>
<connection>
<GID>362</GID>
<name>IN_1</name></connection>
<intersection>-506 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-506,62.5,-505,62.5</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<intersection>-506 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-510.5,78,-506,78</points>
<connection>
<GID>361</GID>
<name>OUT</name></connection>
<intersection>-507.5 4</intersection>
<intersection>-506 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-507.5,75,-507.5,78</points>
<intersection>75 6</intersection>
<intersection>78 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-507.5,75,-505,75</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>-507.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-518.5,79,-518.5,83</points>
<intersection>79 2</intersection>
<intersection>83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-518.5,83,-505,83</points>
<connection>
<GID>362</GID>
<name>IN_0</name></connection>
<intersection>-518.5 0</intersection>
<intersection>-511 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-518.5,79,-516.5,79</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<intersection>-518.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-511,83,-511,94</points>
<intersection>83 1</intersection>
<intersection>94 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-511,94,-496.5,94</points>
<connection>
<GID>352</GID>
<name>OUT</name></connection>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>-511 3</intersection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-518.5,73,-518.5,77</points>
<intersection>73 2</intersection>
<intersection>74 3</intersection>
<intersection>77 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-518.5,77,-516.5,77</points>
<connection>
<GID>361</GID>
<name>IN_1</name></connection>
<intersection>-518.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-518.5,73,-505,73</points>
<connection>
<GID>363</GID>
<name>IN_1</name></connection>
<intersection>-518.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-524,74,-518.5,74</points>
<connection>
<GID>360</GID>
<name>OUT</name></connection>
<intersection>-518.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-533,71,-533,73</points>
<intersection>71 2</intersection>
<intersection>73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-533,73,-530,73</points>
<connection>
<GID>360</GID>
<name>IN_1</name></connection>
<intersection>-533 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-536,71,-533,71</points>
<connection>
<GID>359</GID>
<name>OUT</name></connection>
<intersection>-533 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-533,75,-533,78</points>
<intersection>75 1</intersection>
<intersection>78 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-533,75,-530,75</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>-533 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-536,78,-533,78</points>
<connection>
<GID>358</GID>
<name>OUT</name></connection>
<intersection>-533 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-558.5,70,-542,70</points>
<connection>
<GID>359</GID>
<name>IN_1</name></connection>
<intersection>-558.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-558.5,70,-558.5,72</points>
<intersection>70 1</intersection>
<intersection>71.5 9</intersection>
<intersection>72 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-558.5,72,-556,72</points>
<intersection>-558.5 4</intersection>
<intersection>-556 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-556,72,-556,73.5</points>
<connection>
<GID>357</GID>
<name>IN_1</name></connection>
<intersection>72 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-563,71.5,-558.5,71.5</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<intersection>-558.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-558.5,79,-542,79</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<intersection>-558.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-558.5,76.5,-558.5,79</points>
<intersection>76.5 9</intersection>
<intersection>77 6</intersection>
<intersection>79 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-558.5,77,-556,77</points>
<intersection>-558.5 4</intersection>
<intersection>-556 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-556,75.5,-556,77</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<intersection>77 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-564,76.5,-558.5,76.5</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>-558.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-546,60.5,-546,77</points>
<intersection>60.5 3</intersection>
<intersection>72 6</intersection>
<intersection>74.5 1</intersection>
<intersection>77 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-550,74.5,-546,74.5</points>
<connection>
<GID>357</GID>
<name>OUT</name></connection>
<intersection>-546 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-546,77,-542,77</points>
<connection>
<GID>358</GID>
<name>IN_1</name></connection>
<intersection>-546 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-546,60.5,-505,60.5</points>
<connection>
<GID>365</GID>
<name>IN_1</name></connection>
<intersection>-546 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-546,72,-542,72</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<intersection>-546 0</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-496,74,-496,77</points>
<intersection>74 2</intersection>
<intersection>77 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-496,77,-493,77</points>
<connection>
<GID>364</GID>
<name>IN_1</name></connection>
<intersection>-496 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-499,74,-496,74</points>
<connection>
<GID>363</GID>
<name>OUT</name></connection>
<intersection>-496 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-496,79,-496,82</points>
<intersection>79 1</intersection>
<intersection>82 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-496,79,-493,79</points>
<connection>
<GID>364</GID>
<name>IN_0</name></connection>
<intersection>-496 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-499,82,-496,82</points>
<connection>
<GID>362</GID>
<name>OUT</name></connection>
<intersection>-496 0</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-487,78,-484.5,78</points>
<connection>
<GID>368</GID>
<name>IN_0</name></connection>
<intersection>-487 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-487,78,-487,78</points>
<connection>
<GID>364</GID>
<name>OUT</name></connection>
<intersection>78 1</intersection></vsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-506,29.5,-506,48</points>
<intersection>29.5 2</intersection>
<intersection>45 3</intersection>
<intersection>48 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-506,48,-505,48</points>
<connection>
<GID>375</GID>
<name>IN_1</name></connection>
<intersection>-506 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-506,29.5,-505,29.5</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>-506 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-510.5,45,-506,45</points>
<connection>
<GID>374</GID>
<name>OUT</name></connection>
<intersection>-507.5 4</intersection>
<intersection>-506 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-507.5,42,-507.5,45</points>
<intersection>42 6</intersection>
<intersection>45 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-507.5,42,-505,42</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>-507.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-518.5,46,-518.5,50</points>
<intersection>46 2</intersection>
<intersection>50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-518.5,50,-505,50</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>-518.5 0</intersection>
<intersection>-510 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-518.5,46,-516.5,46</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<intersection>-518.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-510,50,-510,61.5</points>
<intersection>50 1</intersection>
<intersection>61.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-510,61.5,-496,61.5</points>
<connection>
<GID>365</GID>
<name>OUT</name></connection>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<intersection>-510 3</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-518.5,40,-518.5,44</points>
<intersection>40 2</intersection>
<intersection>41 3</intersection>
<intersection>44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-518.5,44,-516.5,44</points>
<connection>
<GID>374</GID>
<name>IN_1</name></connection>
<intersection>-518.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-518.5,40,-505,40</points>
<connection>
<GID>376</GID>
<name>IN_1</name></connection>
<intersection>-518.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-524,41,-518.5,41</points>
<connection>
<GID>373</GID>
<name>OUT</name></connection>
<intersection>-518.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-533,38,-533,40</points>
<intersection>38 2</intersection>
<intersection>40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-533,40,-530,40</points>
<connection>
<GID>373</GID>
<name>IN_1</name></connection>
<intersection>-533 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-536,38,-533,38</points>
<connection>
<GID>372</GID>
<name>OUT</name></connection>
<intersection>-533 0</intersection></hsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-533,42,-533,45</points>
<intersection>42 1</intersection>
<intersection>45 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-533,42,-530,42</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<intersection>-533 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-536,45,-533,45</points>
<connection>
<GID>371</GID>
<name>OUT</name></connection>
<intersection>-533 0</intersection></hsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-558.5,37,-542,37</points>
<connection>
<GID>372</GID>
<name>IN_1</name></connection>
<intersection>-558.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-558.5,37,-558.5,39</points>
<intersection>37 1</intersection>
<intersection>39 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-562.5,39,-556,39</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>-558.5 4</intersection>
<intersection>-556 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-556,39,-556,40.5</points>
<connection>
<GID>370</GID>
<name>IN_1</name></connection>
<intersection>39 6</intersection></vsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-558.5,46,-542,46</points>
<connection>
<GID>371</GID>
<name>IN_0</name></connection>
<intersection>-558.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-558.5,44,-558.5,46</points>
<intersection>44 6</intersection>
<intersection>44.5 9</intersection>
<intersection>46 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-558.5,44,-556,44</points>
<intersection>-558.5 4</intersection>
<intersection>-556 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-556,42.5,-556,44</points>
<connection>
<GID>370</GID>
<name>IN_0</name></connection>
<intersection>44 6</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-563.5,44.5,-558.5,44.5</points>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<intersection>-558.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-546,27.5,-546,44</points>
<intersection>27.5 3</intersection>
<intersection>39 6</intersection>
<intersection>41.5 1</intersection>
<intersection>44 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-550,41.5,-546,41.5</points>
<connection>
<GID>370</GID>
<name>OUT</name></connection>
<intersection>-546 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-546,44,-542,44</points>
<connection>
<GID>371</GID>
<name>IN_1</name></connection>
<intersection>-546 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-546,27.5,-505,27.5</points>
<connection>
<GID>378</GID>
<name>IN_1</name></connection>
<intersection>-546 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-546,39,-542,39</points>
<connection>
<GID>372</GID>
<name>IN_0</name></connection>
<intersection>-546 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-496,41,-496,44</points>
<intersection>41 2</intersection>
<intersection>44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-496,44,-493,44</points>
<connection>
<GID>377</GID>
<name>IN_1</name></connection>
<intersection>-496 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-499,41,-496,41</points>
<connection>
<GID>376</GID>
<name>OUT</name></connection>
<intersection>-496 0</intersection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-496,46,-496,49</points>
<intersection>46 1</intersection>
<intersection>49 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-496,46,-493,46</points>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>-496 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-499,49,-496,49</points>
<connection>
<GID>375</GID>
<name>OUT</name></connection>
<intersection>-496 0</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-487,45,-484.5,45</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>-487 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-487,45,-487,45</points>
<connection>
<GID>377</GID>
<name>OUT</name></connection>
<intersection>45 1</intersection></vsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-499,28.5,-496,28.5</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<intersection>-499 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-499,28.5,-499,28.5</points>
<connection>
<GID>378</GID>
<name>OUT</name></connection>
<intersection>28.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-506.5,125.5,-506.5,144</points>
<intersection>125.5 2</intersection>
<intersection>141 3</intersection>
<intersection>144 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-506.5,144,-505.5,144</points>
<connection>
<GID>286</GID>
<name>IN_1</name></connection>
<intersection>-506.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-506.5,125.5,-505.5,125.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>-506.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-511,141,-506.5,141</points>
<connection>
<GID>285</GID>
<name>OUT</name></connection>
<intersection>-508 4</intersection>
<intersection>-506.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-508,138,-508,141</points>
<intersection>138 6</intersection>
<intersection>141 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-508,138,-505.5,138</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>-508 4</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-519,142,-519,150.5</points>
<intersection>142 2</intersection>
<intersection>146 1</intersection>
<intersection>150.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-519,146,-505.5,146</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>-519 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-519,142,-517,142</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>-519 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-546.5,150.5,-519,150.5</points>
<connection>
<GID>327</GID>
<name>OUT</name></connection>
<intersection>-519 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-519,136,-519,140</points>
<intersection>136 2</intersection>
<intersection>137 3</intersection>
<intersection>140 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-519,140,-517,140</points>
<connection>
<GID>285</GID>
<name>IN_1</name></connection>
<intersection>-519 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-519,136,-505.5,136</points>
<connection>
<GID>287</GID>
<name>IN_1</name></connection>
<intersection>-519 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-524.5,137,-519,137</points>
<connection>
<GID>284</GID>
<name>OUT</name></connection>
<intersection>-519 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-533.5,134,-533.5,136</points>
<intersection>134 2</intersection>
<intersection>136 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-533.5,136,-530.5,136</points>
<connection>
<GID>284</GID>
<name>IN_1</name></connection>
<intersection>-533.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-536.5,134,-533.5,134</points>
<connection>
<GID>283</GID>
<name>OUT</name></connection>
<intersection>-533.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-533.5,138,-533.5,141</points>
<intersection>138 1</intersection>
<intersection>141 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-533.5,138,-530.5,138</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>-533.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-536.5,141,-533.5,141</points>
<connection>
<GID>282</GID>
<name>OUT</name></connection>
<intersection>-533.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-559,133,-542.5,133</points>
<connection>
<GID>283</GID>
<name>IN_1</name></connection>
<intersection>-559 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-559,133,-559,135</points>
<intersection>133 1</intersection>
<intersection>135 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-561.5,135,-556.5,135</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>-559 4</intersection>
<intersection>-556.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-556.5,135,-556.5,136.5</points>
<connection>
<GID>281</GID>
<name>IN_1</name></connection>
<intersection>135 6</intersection></vsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-559,142,-542.5,142</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>-559 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-559,140,-559,142</points>
<intersection>140 6</intersection>
<intersection>142 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-562.5,140,-556.5,140</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>-559 4</intersection>
<intersection>-556.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-556.5,138.5,-556.5,140</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>140 6</intersection></vsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-546.5,123.5,-546.5,140</points>
<intersection>123.5 3</intersection>
<intersection>135 6</intersection>
<intersection>137.5 1</intersection>
<intersection>140 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-550.5,137.5,-546.5,137.5</points>
<connection>
<GID>281</GID>
<name>OUT</name></connection>
<intersection>-546.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-546.5,140,-542.5,140</points>
<connection>
<GID>282</GID>
<name>IN_1</name></connection>
<intersection>-546.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-546.5,123.5,-505.5,123.5</points>
<connection>
<GID>289</GID>
<name>IN_1</name></connection>
<intersection>-546.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-546.5,135,-542.5,135</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>-546.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-496.5,137,-496.5,140</points>
<intersection>137 2</intersection>
<intersection>140 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-496.5,140,-493.5,140</points>
<connection>
<GID>288</GID>
<name>IN_1</name></connection>
<intersection>-496.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-499.5,137,-496.5,137</points>
<connection>
<GID>287</GID>
<name>OUT</name></connection>
<intersection>-496.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-496.5,142,-496.5,145</points>
<intersection>142 1</intersection>
<intersection>145 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-496.5,142,-493.5,142</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>-496.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-499.5,145,-496.5,145</points>
<connection>
<GID>286</GID>
<name>OUT</name></connection>
<intersection>-496.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-571,148.5,-571,158.5</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>148.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-571,148.5,-564.5,148.5</points>
<connection>
<GID>325</GID>
<name>IN_1</name></connection>
<intersection>-571 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-567.5,150.5,-567.5,158.5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>150.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-567.5,150.5,-564.5,150.5</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>-567.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-558.5,149.5,-552.5,149.5</points>
<connection>
<GID>325</GID>
<name>OUT</name></connection>
<connection>
<GID>327</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-556,151.5,-556,158.5</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>151.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-556,151.5,-552.5,151.5</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>-556 0</intersection></hsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-487.5,141,-485,141</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>-487.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-487.5,141,-487.5,141</points>
<connection>
<GID>288</GID>
<name>OUT</name></connection>
<intersection>141 1</intersection></vsegment></shape></wire></page 3>
<page 4>
<PageViewport>54.724,-51.8764,108.892,-112.795</PageViewport></page 4>
<page 5>
<PageViewport>-53.2278,36.0834,43.0722,-72.2167</PageViewport></page 5>
<page 6>
<PageViewport>-6.2,4.85,90.1,-103.45</PageViewport></page 6>
<page 7>
<PageViewport>-6.2,4.85,90.1,-103.45</PageViewport></page 7>
<page 8>
<PageViewport>-6.2,4.85,90.1,-103.45</PageViewport></page 8>
<page 9>
<PageViewport>-6.2,4.85,90.1,-103.45</PageViewport></page 9></circuit>