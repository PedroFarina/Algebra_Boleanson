<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-94.4376,85.825,33.9624,-58.575</PageViewport>
<gate>
<ID>198</ID>
<type>AA_TOGGLE</type>
<position>-50,13</position>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>-85.5,13</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>DE_TO</type>
<position>-82.5,24.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>-98,13</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>203</ID>
<type>DE_TO</type>
<position>-47,24.5</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S 2</lparam></gate>
<gate>
<ID>11</ID>
<type>DE_TO</type>
<position>-95,24.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>-36.5,13</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>DE_TO</type>
<position>-33.5,24.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S 3</lparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>-24,13</position>
<input>
<ID>N_in3</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>212</ID>
<type>DE_TO</type>
<position>-18,24.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Output 1</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>0,13</position>
<input>
<ID>N_in3</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>DE_TO</type>
<position>6,24.5</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Output 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>-74,13</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>37</ID>
<type>DE_TO</type>
<position>-71,24.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cin</lparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>25,13</position>
<input>
<ID>N_in3</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>DE_TO</type>
<position>31,24.5</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cout</lparam></gate>
<gate>
<ID>164</ID>
<type>AA_TOGGLE</type>
<position>-62.5,13</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>185</ID>
<type>DE_TO</type>
<position>-59.5,24.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S 1</lparam></gate>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-98,15,-98,24.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-98,24.5,-97,24.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>-98 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-85.5,15,-85.5,24.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-85.5,24.5,-84.5,24.5</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>-85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24,14,-24,24.5</points>
<connection>
<GID>19</GID>
<name>N_in3</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,24.5,-20,24.5</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>-24 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,15,-36.5,24.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,24.5,-35.5,24.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,14,0,24.5</points>
<connection>
<GID>34</GID>
<name>N_in3</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,24.5,4,24.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>0 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74,15,-74,24.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-74,24.5,-73,24.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>-74 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,14,25,24.5</points>
<connection>
<GID>38</GID>
<name>N_in3</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,24.5,29,24.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62.5,15,-62.5,24.5</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62.5,24.5,-61.5,24.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>-62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-50,15,-50,24.5</points>
<connection>
<GID>198</GID>
<name>OUT_0</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-50,24.5,-49,24.5</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>-50 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-106.35,82.5296,164.494,-222.064</PageViewport>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>14.5,-19</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_OR2</type>
<position>14.5,-25</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AI_XOR2</type>
<position>14.5,-31</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>DA_FROM</type>
<position>35,-10.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S 1</lparam></gate>
<gate>
<ID>17</ID>
<type>DA_FROM</type>
<position>39.5,-10.5</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S 2</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>43.5,-10.5</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID S 3</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_AND2</type>
<position>14.5,-105.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>BA_NAND2</type>
<position>14.5,-37.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_OR2</type>
<position>14.5,-111.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>BE_NOR2</type>
<position>14.5,-44</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AI_XOR2</type>
<position>14.5,-117.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AO_XNOR2</type>
<position>14.5,-50.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>BA_NAND2</type>
<position>14.5,-124</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>AI_MUX_8x1</type>
<position>39.5,-32.5</position>
<input>
<ID>IN_1</ID>37 </input>
<input>
<ID>IN_2</ID>13 </input>
<input>
<ID>IN_3</ID>12 </input>
<input>
<ID>IN_4</ID>11 </input>
<input>
<ID>IN_5</ID>10 </input>
<input>
<ID>IN_6</ID>9 </input>
<input>
<ID>IN_7</ID>8 </input>
<output>
<ID>OUT</ID>14 </output>
<input>
<ID>SEL_0</ID>19 </input>
<input>
<ID>SEL_1</ID>18 </input>
<input>
<ID>SEL_2</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>28</ID>
<type>BE_NOR2</type>
<position>14.5,-130.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>AO_XNOR2</type>
<position>14.5,-137</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AI_MUX_8x1</type>
<position>39.5,-119</position>
<input>
<ID>IN_1</ID>44 </input>
<input>
<ID>IN_2</ID>27 </input>
<input>
<ID>IN_3</ID>26 </input>
<input>
<ID>IN_4</ID>25 </input>
<input>
<ID>IN_5</ID>24 </input>
<input>
<ID>IN_6</ID>23 </input>
<input>
<ID>IN_7</ID>22 </input>
<output>
<ID>OUT</ID>28 </output>
<input>
<ID>SEL_0</ID>19 </input>
<input>
<ID>SEL_1</ID>18 </input>
<input>
<ID>SEL_2</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>31</ID>
<type>DA_FROM</type>
<position>-16,-96</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>32</ID>
<type>DA_FROM</type>
<position>-11,-96</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>33</ID>
<type>DE_TO</type>
<position>55.5,-105</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Output 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AI_XOR2</type>
<position>-5,-59.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_AND2</type>
<position>-5,-69</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AI_XOR2</type>
<position>14,-58.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_AND2</type>
<position>14,-65</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>DA_FROM</type>
<position>3,-12.5</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID Cin</lparam></gate>
<gate>
<ID>45</ID>
<type>AE_OR2</type>
<position>26.5,-68</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AI_XOR2</type>
<position>-5,-145.5</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_AND2</type>
<position>-5,-155</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>AI_XOR2</type>
<position>14,-144.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_AND2</type>
<position>14,-151</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>AE_OR2</type>
<position>26.5,-154</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>DE_TO</type>
<position>52,-154</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID Cout</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>17.5,12.5</position>
<gparam>LABEL_TEXT Unidade L�gica Aritim�tica</gparam>
<gparam>TEXT_HEIGHT 6</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>DA_FROM</type>
<position>-16,-10.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>90</ID>
<type>DA_FROM</type>
<position>-11,-10.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>145</ID>
<type>DE_TO</type>
<position>55.5,-17.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID Output 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-70,-11,-12.5</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>-70 15</intersection>
<intersection>-58.5 13</intersection>
<intersection>-49.5 11</intersection>
<intersection>-43 8</intersection>
<intersection>-36.5 9</intersection>
<intersection>-30 4</intersection>
<intersection>-24 5</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11,-18,11.5,-18</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-11,-30,11.5,-30</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-11,-24,11.5,-24</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-11,-43,11.5,-43</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-11,-36.5,11.5,-36.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-11,-49.5,11.5,-49.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-11,-58.5,-8,-58.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-11,-70,-8,-70</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>-11 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-68,-16,-12.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>-68 15</intersection>
<intersection>-60.5 13</intersection>
<intersection>-51.5 10</intersection>
<intersection>-45 11</intersection>
<intersection>-38.5 7</intersection>
<intersection>-32 4</intersection>
<intersection>-26 5</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-20,11.5,-20</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-16,-32,11.5,-32</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-16,-26,11.5,-26</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-16,-38.5,11.5,-38.5</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-16,-51.5,11.5,-51.5</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-16,-45,11.5,-45</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-16,-60.5,-8,-60.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-16,-68,-8,-68</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-29,25.5,-19</points>
<intersection>-29 1</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-29,36.5,-29</points>
<connection>
<GID>27</GID>
<name>IN_7</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-19,25.5,-19</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-30,25,-25</points>
<intersection>-30 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-30,36.5,-30</points>
<connection>
<GID>27</GID>
<name>IN_6</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-25,25,-25</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-31,36.5,-31</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<connection>
<GID>27</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-37.5,24,-32</points>
<intersection>-37.5 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-32,36.5,-32</points>
<connection>
<GID>27</GID>
<name>IN_4</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-37.5,24,-37.5</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-44,24.5,-33</points>
<intersection>-44 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-33,36.5,-33</points>
<connection>
<GID>27</GID>
<name>IN_3</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-44,24.5,-44</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-50.5,25,-34</points>
<intersection>-50.5 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-34,36.5,-34</points>
<connection>
<GID>27</GID>
<name>IN_2</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-50.5,25,-50.5</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-32.5,55.5,-19.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-32.5,55.5,-32.5</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-113.5,38.5,-19.5</points>
<connection>
<GID>27</GID>
<name>SEL_2</name></connection>
<connection>
<GID>30</GID>
<name>SEL_2</name></connection>
<intersection>-19.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>35,-19.5,35,-12.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35,-19.5,38.5,-19.5</points>
<intersection>35 1</intersection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-113.5,39.5,-12.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>SEL_1</name></connection>
<connection>
<GID>30</GID>
<name>SEL_1</name></connection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-113.5,40.5,-19.5</points>
<connection>
<GID>27</GID>
<name>SEL_0</name></connection>
<connection>
<GID>30</GID>
<name>SEL_0</name></connection>
<intersection>-19.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>43.5,-19.5,43.5,-12.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>40.5,-19.5,43.5,-19.5</points>
<intersection>40.5 0</intersection>
<intersection>43.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11,-156,-11,-98</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>-156 28</intersection>
<intersection>-144.5 26</intersection>
<intersection>-136 11</intersection>
<intersection>-129.5 8</intersection>
<intersection>-123 9</intersection>
<intersection>-116.5 4</intersection>
<intersection>-110.5 5</intersection>
<intersection>-104.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-11,-104.5,11.5,-104.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-11,-116.5,11.5,-116.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-11,-110.5,11.5,-110.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-11,-129.5,11.5,-129.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-11,-123,11.5,-123</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-11,-136,11.5,-136</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>-11,-144.5,-8,-144.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>-11 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-11,-156,-8,-156</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>-11 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-115.5,25.5,-105.5</points>
<intersection>-115.5 1</intersection>
<intersection>-105.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-115.5,36.5,-115.5</points>
<connection>
<GID>30</GID>
<name>IN_7</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-105.5,25.5,-105.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-116.5,25,-111.5</points>
<intersection>-116.5 1</intersection>
<intersection>-111.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-116.5,36.5,-116.5</points>
<connection>
<GID>30</GID>
<name>IN_6</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-111.5,25,-111.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-117.5,36.5,-117.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<connection>
<GID>30</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-124,24,-118.5</points>
<intersection>-124 2</intersection>
<intersection>-118.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-118.5,36.5,-118.5</points>
<connection>
<GID>30</GID>
<name>IN_4</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-124,24,-124</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-130.5,24.5,-119.5</points>
<intersection>-130.5 2</intersection>
<intersection>-119.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-119.5,36.5,-119.5</points>
<connection>
<GID>30</GID>
<name>IN_3</name></connection>
<intersection>24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-130.5,24.5,-130.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-137,25,-120.5</points>
<intersection>-137 2</intersection>
<intersection>-120.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-120.5,36.5,-120.5</points>
<connection>
<GID>30</GID>
<name>IN_2</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-137,25,-137</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-119,55.5,-107</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>-119 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-119,55.5,-119</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-59.5,11,-59.5</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>8.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>8.5,-64,8.5,-59.5</points>
<intersection>-64 4</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>8.5,-64,11,-64</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>8.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-66,3,-14.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-66 3</intersection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,-57.5,11,-57.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>3,-66,11,-66</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-67,20,-65</points>
<intersection>-67 2</intersection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-65,20,-65</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20,-67,23.5,-67</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-69,23.5,-69</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<connection>
<GID>45</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-58.5,26.5,-35</points>
<intersection>-58.5 2</intersection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-35,36.5,-35</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-58.5,26.5,-58.5</points>
<connection>
<GID>42</GID>
<name>OUT</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-154,-16,-98</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-154 15</intersection>
<intersection>-146.5 13</intersection>
<intersection>-138 27</intersection>
<intersection>-131.5 28</intersection>
<intersection>-125 24</intersection>
<intersection>-118.5 21</intersection>
<intersection>-112.5 22</intersection>
<intersection>-106.5 18</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-16,-146.5,-8,-146.5</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-16,-154,-8,-154</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>18</ID>
<points>-16,-106.5,11.5,-106.5</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>-16,-118.5,11.5,-118.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>-16,-112.5,11.5,-112.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>-16,-125,11.5,-125</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>-16,-138,11.5,-138</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>-16,-131.5,11.5,-131.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-145.5,11,-145.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>8.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>8.5,-150,8.5,-145.5</points>
<intersection>-150 4</intersection>
<intersection>-145.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>8.5,-150,11,-150</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>8.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-152,3,-82.5</points>
<intersection>-152 3</intersection>
<intersection>-143.5 1</intersection>
<intersection>-82.5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,-143.5,11,-143.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>3,-152,11,-152</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>3,-82.5,32.5,-82.5</points>
<intersection>3 0</intersection>
<intersection>32.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>32.5,-82.5,32.5,-68</points>
<intersection>-82.5 5</intersection>
<intersection>-68 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>29.5,-68,32.5,-68</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>32.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-153,20,-151</points>
<intersection>-153 2</intersection>
<intersection>-151 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-151,20,-151</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20,-153,23.5,-153</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2,-155,23.5,-155</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<connection>
<GID>51</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-144.5,26.5,-121.5</points>
<intersection>-144.5 2</intersection>
<intersection>-121.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-121.5,36.5,-121.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-144.5,26.5,-144.5</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-154,50,-154</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>29.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>29.5,-154,29.5,-154</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>-154 1</intersection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>-18.6403,14.5271,77.6597,-93.7729</PageViewport></page 2>
<page 3>
<PageViewport>-635.271,212.555,-364.426,-92.0405</PageViewport></page 3>
<page 4>
<PageViewport>54.7234,-51.8764,108.892,-112.795</PageViewport></page 4>
<page 5>
<PageViewport>-53.2278,36.0834,43.0722,-72.2167</PageViewport></page 5>
<page 6>
<PageViewport>-6.2,4.85,90.1,-103.45</PageViewport></page 6>
<page 7>
<PageViewport>-6.2,4.85,90.1,-103.45</PageViewport></page 7>
<page 8>
<PageViewport>-6.2,4.85,90.1,-103.45</PageViewport></page 8>
<page 9>
<PageViewport>-6.2,4.85,90.1,-103.45</PageViewport></page 9></circuit>