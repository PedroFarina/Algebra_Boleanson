<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-100.146,116.2,28.2536,-28.2</PageViewport>
<gate>
<ID>198</ID>
<type>AA_TOGGLE</type>
<position>-38.5,13</position>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>203</ID>
<type>DE_TO</type>
<position>-35.5,24.5</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>212</ID>
<type>DE_TO</type>
<position>-18,24.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S</lparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>-24,13</position>
<input>
<ID>N_in3</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>AA_TOGGLE</type>
<position>-51,13</position>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>185</ID>
<type>DE_TO</type>
<position>-48,24.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24,14,-24,24.5</points>
<connection>
<GID>19</GID>
<name>N_in3</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,24.5,-20,24.5</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>-24 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51,15,-51,24.5</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-51,24.5,-50,24.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>-51 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-38.5,15,-38.5,24.5</points>
<connection>
<GID>198</GID>
<name>OUT_0</name></connection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-38.5,24.5,-37.5,24.5</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>-38.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-27.0037,9.81466,58.6932,-86.561</PageViewport>
<gate>
<ID>4</ID>
<type>AA_AND2</type>
<position>14.5,-19</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_OR2</type>
<position>14.5,-25</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AI_XOR2</type>
<position>14.5,-31</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>BA_NAND2</type>
<position>14.5,-37.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>BE_NOR2</type>
<position>14.5,-44</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AO_XNOR2</type>
<position>14.5,-50.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>AI_MUX_8x1</type>
<position>39.5,-32.5</position>
<input>
<ID>IN_2</ID>13 </input>
<input>
<ID>IN_3</ID>12 </input>
<input>
<ID>IN_4</ID>11 </input>
<input>
<ID>IN_5</ID>10 </input>
<input>
<ID>IN_6</ID>9 </input>
<input>
<ID>IN_7</ID>8 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>89</ID>
<type>DA_FROM</type>
<position>-16,-10.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>90</ID>
<type>DA_FROM</type>
<position>3,-11</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 270</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>145</ID>
<type>DE_TO</type>
<position>48,-20</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID S</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-49.5,3,-13</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>-49.5 11</intersection>
<intersection>-43 8</intersection>
<intersection>-36.5 9</intersection>
<intersection>-30 4</intersection>
<intersection>-24 5</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,-18,11.5,-18</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>3,-30,11.5,-30</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>3,-24,11.5,-24</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>3,-43,11.5,-43</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>3,-36.5,11.5,-36.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>3,-49.5,11.5,-49.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-16,-51.5,-16,-12.5</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>-51.5 10</intersection>
<intersection>-45 11</intersection>
<intersection>-38.5 7</intersection>
<intersection>-32 4</intersection>
<intersection>-26 5</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-16,-20,11.5,-20</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-16,-32,11.5,-32</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-16,-26,11.5,-26</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-16,-38.5,11.5,-38.5</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>-16,-51.5,11.5,-51.5</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-16,-45,11.5,-45</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>-16 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-29,25,-19</points>
<intersection>-29 1</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-29,36.5,-29</points>
<connection>
<GID>27</GID>
<name>IN_7</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-19,25,-19</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-30,25,-25</points>
<intersection>-30 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-30,36.5,-30</points>
<connection>
<GID>27</GID>
<name>IN_6</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-25,25,-25</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-31,36.5,-31</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<connection>
<GID>27</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-37.5,25,-32</points>
<intersection>-37.5 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-32,36.5,-32</points>
<connection>
<GID>27</GID>
<name>IN_4</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-37.5,25,-37.5</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-44,25,-33</points>
<intersection>-44 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-33,36.5,-33</points>
<connection>
<GID>27</GID>
<name>IN_3</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-44,25,-44</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-50.5,25,-34</points>
<intersection>-50.5 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-34,36.5,-34</points>
<connection>
<GID>27</GID>
<name>IN_2</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-50.5,25,-50.5</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-32.5,48,-22</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-32.5,48,-32.5</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-18.6403,14.5271,77.6597,-93.7729</PageViewport></page 2>
<page 3>
<PageViewport>-635.271,212.555,-364.426,-92.0405</PageViewport></page 3>
<page 4>
<PageViewport>54.7235,-51.8764,108.892,-112.795</PageViewport></page 4>
<page 5>
<PageViewport>-53.2278,36.0834,43.0722,-72.2167</PageViewport></page 5>
<page 6>
<PageViewport>-6.2,4.85,90.1,-103.45</PageViewport></page 6>
<page 7>
<PageViewport>-6.2,4.85,90.1,-103.45</PageViewport></page 7>
<page 8>
<PageViewport>-6.2,4.85,90.1,-103.45</PageViewport></page 8>
<page 9>
<PageViewport>-6.2,4.85,90.1,-103.45</PageViewport></page 9></circuit>