<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-35.887,1.44764,116.531,-78.0191</PageViewport>
<gate>
<ID>2</ID>
<type>DA_FROM</type>
<position>14.5,-10.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DME0</lparam></gate>
<gate>
<ID>3</ID>
<type>DA_FROM</type>
<position>14.5,-13.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DME1</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_SMALL_INVERTER</type>
<position>36.5,-21</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AE_SMALL_INVERTER</type>
<position>40.5,-21</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_AND3</type>
<position>50,-40.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>2 </input>
<input>
<ID>IN_2</ID>7 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_AND3</type>
<position>50,-51</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>1 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND3</type>
<position>50,-30.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>7 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_AND3</type>
<position>50.5,-60.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<input>
<ID>IN_2</ID>7 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>13</ID>
<type>DA_FROM</type>
<position>6,-37</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DMI</lparam></gate>
<gate>
<ID>15</ID>
<type>DE_TO</type>
<position>56.5,-30.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DM0</lparam></gate>
<gate>
<ID>16</ID>
<type>DE_TO</type>
<position>57,-40.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DM1</lparam></gate>
<gate>
<ID>17</ID>
<type>DE_TO</type>
<position>57,-51</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DM2</lparam></gate>
<gate>
<ID>18</ID>
<type>DE_TO</type>
<position>57.5,-60.5</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DM3</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-60.5,23,-13.5</points>
<intersection>-60.5 2</intersection>
<intersection>-53 5</intersection>
<intersection>-19 3</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-13.5,23,-13.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-60.5,47.5,-60.5</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>23,-19,40.5,-19</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>23,-53,47,-53</points>
<connection>
<GID>9</GID>
<name>IN_2</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-58.5,26.5,-10.5</points>
<intersection>-58.5 5</intersection>
<intersection>-40.5 2</intersection>
<intersection>-19 3</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-10.5,26.5,-10.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-40.5,47,-40.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26.5,-19,36.5,-19</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>26.5,-58.5,47.5,-58.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-38.5,40.5,-23</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>-38.5 3</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-28.5,47,-28.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>40.5,-38.5,47,-38.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-51,36.5,-23</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>-51 3</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-30.5,47,-30.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36.5,-51,47,-51</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8,-37,16,-37</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>16 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16,-62.5,16,-32.5</points>
<intersection>-62.5 5</intersection>
<intersection>-49 6</intersection>
<intersection>-42.5 7</intersection>
<intersection>-37 1</intersection>
<intersection>-32.5 10</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>16,-62.5,47.5,-62.5</points>
<connection>
<GID>11</GID>
<name>IN_2</name></connection>
<intersection>16 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>16,-49,47,-49</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>16 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>16,-42.5,47,-42.5</points>
<connection>
<GID>8</GID>
<name>IN_2</name></connection>
<intersection>16 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>16,-32.5,47,-32.5</points>
<connection>
<GID>10</GID>
<name>IN_2</name></connection>
<intersection>16 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-40.5,55,-40.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-30.5,54.5,-30.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53,-51,55,-51</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<connection>
<GID>17</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>53.5,-60.5,55.5,-60.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<connection>
<GID>11</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-63.5514,6.7459,106.939,-82.143</PageViewport>
<gate>
<ID>20</ID>
<type>DA_FROM</type>
<position>10,-5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ME0</lparam></gate>
<gate>
<ID>21</ID>
<type>DA_FROM</type>
<position>10,-8</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ME1</lparam></gate>
<gate>
<ID>23</ID>
<type>AE_MUX_4x1</type>
<position>23,-17.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>15 </input>
<input>
<ID>IN_3</ID>14 </input>
<output>
<ID>OUT</ID>30 </output>
<input>
<ID>SEL_0</ID>13 </input>
<input>
<ID>SEL_1</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>25</ID>
<type>DA_FROM</type>
<position>3.5,-14.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MD0</lparam></gate>
<gate>
<ID>26</ID>
<type>DA_FROM</type>
<position>3.5,-16.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MC0</lparam></gate>
<gate>
<ID>27</ID>
<type>DA_FROM</type>
<position>3.5,-18.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MB0</lparam></gate>
<gate>
<ID>28</ID>
<type>DA_FROM</type>
<position>3.5,-20.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MA0</lparam></gate>
<gate>
<ID>29</ID>
<type>AE_MUX_4x1</type>
<position>23,-34</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>20 </input>
<input>
<ID>IN_2</ID>19 </input>
<input>
<ID>IN_3</ID>18 </input>
<output>
<ID>OUT</ID>31 </output>
<input>
<ID>SEL_0</ID>13 </input>
<input>
<ID>SEL_1</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>30</ID>
<type>AE_MUX_4x1</type>
<position>23,-49.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>24 </input>
<input>
<ID>IN_2</ID>23 </input>
<input>
<ID>IN_3</ID>22 </input>
<output>
<ID>OUT</ID>32 </output>
<input>
<ID>SEL_0</ID>13 </input>
<input>
<ID>SEL_1</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_MUX_4x1</type>
<position>23,-65.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>28 </input>
<input>
<ID>IN_2</ID>27 </input>
<input>
<ID>IN_3</ID>26 </input>
<output>
<ID>OUT</ID>33 </output>
<input>
<ID>SEL_0</ID>13 </input>
<input>
<ID>SEL_1</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>32</ID>
<type>DA_FROM</type>
<position>3.5,-31</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MD1</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>3.5,-33</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MC1</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>3.5,-35</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MB1</lparam></gate>
<gate>
<ID>35</ID>
<type>DA_FROM</type>
<position>3.5,-37</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MA1</lparam></gate>
<gate>
<ID>36</ID>
<type>DA_FROM</type>
<position>2.5,-46.5</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MD2</lparam></gate>
<gate>
<ID>37</ID>
<type>DA_FROM</type>
<position>2.5,-48.5</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MC2</lparam></gate>
<gate>
<ID>38</ID>
<type>DA_FROM</type>
<position>2.5,-50.5</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MB2</lparam></gate>
<gate>
<ID>39</ID>
<type>DA_FROM</type>
<position>2.5,-52.5</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MA2</lparam></gate>
<gate>
<ID>40</ID>
<type>DA_FROM</type>
<position>2.5,-62</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MD3</lparam></gate>
<gate>
<ID>41</ID>
<type>DA_FROM</type>
<position>2.5,-64</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MC3</lparam></gate>
<gate>
<ID>42</ID>
<type>DA_FROM</type>
<position>2.5,-66</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MB3</lparam></gate>
<gate>
<ID>43</ID>
<type>DA_FROM</type>
<position>2.5,-68</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MA3</lparam></gate>
<gate>
<ID>45</ID>
<type>DE_TO</type>
<position>30,-17.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M0</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>29.5,-34</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M1</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>29.5,-49.5</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M2</lparam></gate>
<gate>
<ID>48</ID>
<type>DE_TO</type>
<position>29.5,-65.5</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M3</lparam></gate>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-60.5,23,-8</points>
<connection>
<GID>31</GID>
<name>SEL_1</name></connection>
<connection>
<GID>30</GID>
<name>SEL_1</name></connection>
<connection>
<GID>23</GID>
<name>SEL_1</name></connection>
<connection>
<GID>29</GID>
<name>SEL_1</name></connection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-8,23,-8</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-60.5,24,-5</points>
<connection>
<GID>31</GID>
<name>SEL_0</name></connection>
<connection>
<GID>30</GID>
<name>SEL_0</name></connection>
<connection>
<GID>23</GID>
<name>SEL_0</name></connection>
<connection>
<GID>29</GID>
<name>SEL_0</name></connection>
<intersection>-5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-5,24,-5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,-14.5,20,-14.5</points>
<connection>
<GID>23</GID>
<name>IN_3</name></connection>
<connection>
<GID>25</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,-16.5,20,-16.5</points>
<connection>
<GID>23</GID>
<name>IN_2</name></connection>
<connection>
<GID>26</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,-18.5,20,-18.5</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<connection>
<GID>27</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,-20.5,20,-20.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,-31,20,-31</points>
<connection>
<GID>29</GID>
<name>IN_3</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,-33,20,-33</points>
<connection>
<GID>29</GID>
<name>IN_2</name></connection>
<connection>
<GID>33</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,-35,20,-35</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<connection>
<GID>34</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>5.5,-37,20,-37</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<connection>
<GID>35</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-46.5,20,-46.5</points>
<connection>
<GID>30</GID>
<name>IN_3</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-48.5,20,-48.5</points>
<connection>
<GID>30</GID>
<name>IN_2</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-50.5,20,-50.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-52.5,20,-52.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-62,20,-62</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>20 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20,-62.5,20,-62</points>
<connection>
<GID>31</GID>
<name>IN_3</name></connection>
<intersection>-62 1</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-64,20,-64</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>20 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20,-64.5,20,-64</points>
<connection>
<GID>31</GID>
<name>IN_2</name></connection>
<intersection>-64 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-66,20,-66</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>20 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20,-66.5,20,-66</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>-66 1</intersection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4.5,-68,20,-68</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>20 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20,-68.5,20,-68</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-68 1</intersection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-17.5,28,-17.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<connection>
<GID>23</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-34,27.5,-34</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<connection>
<GID>29</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-49.5,27.5,-49.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<connection>
<GID>30</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-65.5,27.5,-65.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<connection>
<GID>48</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-83.0916,-16.1006,187.875,-157.375</PageViewport>
<gate>
<ID>50</ID>
<type>AE_DFF_LOW_NT</type>
<position>13.5,-23</position>
<input>
<ID>IN_0</ID>35 </input>
<output>
<ID>OUT_0</ID>42 </output>
<input>
<ID>clock</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>51</ID>
<type>AE_DFF_LOW_NT</type>
<position>24,-23</position>
<input>
<ID>IN_0</ID>36 </input>
<output>
<ID>OUT_0</ID>41 </output>
<input>
<ID>clock</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>52</ID>
<type>AE_DFF_LOW_NT</type>
<position>34,-23</position>
<input>
<ID>IN_0</ID>37 </input>
<output>
<ID>OUT_0</ID>40 </output>
<input>
<ID>clock</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>53</ID>
<type>AE_DFF_LOW_NT</type>
<position>43,-23</position>
<input>
<ID>IN_0</ID>38 </input>
<output>
<ID>OUT_0</ID>39 </output>
<input>
<ID>clock</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>55</ID>
<type>DA_FROM</type>
<position>0,-31.5</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DM0</lparam></gate>
<gate>
<ID>57</ID>
<type>DA_FROM</type>
<position>1,-37.5</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In3</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>1,-40.5</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In2</lparam></gate>
<gate>
<ID>59</ID>
<type>DA_FROM</type>
<position>1,-43.5</position>
<input>
<ID>IN_0</ID>37 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In1</lparam></gate>
<gate>
<ID>60</ID>
<type>DA_FROM</type>
<position>1,-46.5</position>
<input>
<ID>IN_0</ID>38 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In0</lparam></gate>
<gate>
<ID>64</ID>
<type>DE_TO</type>
<position>50,-7.5</position>
<input>
<ID>IN_0</ID>42 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MA3</lparam></gate>
<gate>
<ID>65</ID>
<type>DE_TO</type>
<position>50,-10.5</position>
<input>
<ID>IN_0</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MA2</lparam></gate>
<gate>
<ID>66</ID>
<type>DE_TO</type>
<position>50,-13.5</position>
<input>
<ID>IN_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MA1</lparam></gate>
<gate>
<ID>67</ID>
<type>DE_TO</type>
<position>50,-17</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MA0</lparam></gate>
<gate>
<ID>68</ID>
<type>AE_DFF_LOW_NT</type>
<position>9,-69.5</position>
<input>
<ID>IN_0</ID>44 </input>
<output>
<ID>OUT_0</ID>51 </output>
<input>
<ID>clock</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>69</ID>
<type>AE_DFF_LOW_NT</type>
<position>19.5,-69.5</position>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>50 </output>
<input>
<ID>clock</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>70</ID>
<type>AE_DFF_LOW_NT</type>
<position>29.5,-69.5</position>
<input>
<ID>IN_0</ID>46 </input>
<output>
<ID>OUT_0</ID>49 </output>
<input>
<ID>clock</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_DFF_LOW_NT</type>
<position>38.5,-69.5</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>48 </output>
<input>
<ID>clock</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>72</ID>
<type>DA_FROM</type>
<position>-4.5,-78</position>
<input>
<ID>IN_0</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DM1</lparam></gate>
<gate>
<ID>73</ID>
<type>DA_FROM</type>
<position>-3.5,-84</position>
<input>
<ID>IN_0</ID>44 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In3</lparam></gate>
<gate>
<ID>74</ID>
<type>DA_FROM</type>
<position>-3.5,-87</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In2</lparam></gate>
<gate>
<ID>75</ID>
<type>DA_FROM</type>
<position>-3.5,-90</position>
<input>
<ID>IN_0</ID>46 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In1</lparam></gate>
<gate>
<ID>76</ID>
<type>DA_FROM</type>
<position>-3.5,-93</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In0</lparam></gate>
<gate>
<ID>77</ID>
<type>DE_TO</type>
<position>45.5,-54</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MB3</lparam></gate>
<gate>
<ID>78</ID>
<type>DE_TO</type>
<position>45.5,-57</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MB2</lparam></gate>
<gate>
<ID>79</ID>
<type>DE_TO</type>
<position>45.5,-60</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MB1</lparam></gate>
<gate>
<ID>80</ID>
<type>DE_TO</type>
<position>45.5,-63.5</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MB0</lparam></gate>
<gate>
<ID>81</ID>
<type>AE_DFF_LOW_NT</type>
<position>14,-114.5</position>
<input>
<ID>IN_0</ID>53 </input>
<output>
<ID>OUT_0</ID>60 </output>
<input>
<ID>clock</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>82</ID>
<type>AE_DFF_LOW_NT</type>
<position>24.5,-114.5</position>
<input>
<ID>IN_0</ID>54 </input>
<output>
<ID>OUT_0</ID>59 </output>
<input>
<ID>clock</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>83</ID>
<type>AE_DFF_LOW_NT</type>
<position>34.5,-114.5</position>
<input>
<ID>IN_0</ID>55 </input>
<output>
<ID>OUT_0</ID>58 </output>
<input>
<ID>clock</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>84</ID>
<type>AE_DFF_LOW_NT</type>
<position>43.5,-114.5</position>
<input>
<ID>IN_0</ID>56 </input>
<output>
<ID>OUT_0</ID>57 </output>
<input>
<ID>clock</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>85</ID>
<type>DA_FROM</type>
<position>0.5,-123</position>
<input>
<ID>IN_0</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DM2</lparam></gate>
<gate>
<ID>86</ID>
<type>DA_FROM</type>
<position>1.5,-129</position>
<input>
<ID>IN_0</ID>53 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In3</lparam></gate>
<gate>
<ID>87</ID>
<type>DA_FROM</type>
<position>1.5,-132</position>
<input>
<ID>IN_0</ID>54 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In2</lparam></gate>
<gate>
<ID>88</ID>
<type>DA_FROM</type>
<position>1.5,-135</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In1</lparam></gate>
<gate>
<ID>89</ID>
<type>DA_FROM</type>
<position>1.5,-138</position>
<input>
<ID>IN_0</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In0</lparam></gate>
<gate>
<ID>90</ID>
<type>DE_TO</type>
<position>50.5,-99</position>
<input>
<ID>IN_0</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MC3</lparam></gate>
<gate>
<ID>91</ID>
<type>DE_TO</type>
<position>50.5,-102</position>
<input>
<ID>IN_0</ID>59 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MC2</lparam></gate>
<gate>
<ID>92</ID>
<type>DE_TO</type>
<position>50.5,-105</position>
<input>
<ID>IN_0</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MC1</lparam></gate>
<gate>
<ID>93</ID>
<type>DE_TO</type>
<position>50.5,-108.5</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MC0</lparam></gate>
<gate>
<ID>94</ID>
<type>AE_DFF_LOW_NT</type>
<position>87,-60.5</position>
<input>
<ID>IN_0</ID>62 </input>
<output>
<ID>OUT_0</ID>69 </output>
<input>
<ID>clock</ID>61 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>95</ID>
<type>AE_DFF_LOW_NT</type>
<position>97.5,-60.5</position>
<input>
<ID>IN_0</ID>63 </input>
<output>
<ID>OUT_0</ID>68 </output>
<input>
<ID>clock</ID>61 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>96</ID>
<type>AE_DFF_LOW_NT</type>
<position>107.5,-60.5</position>
<input>
<ID>IN_0</ID>64 </input>
<output>
<ID>OUT_0</ID>67 </output>
<input>
<ID>clock</ID>61 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>97</ID>
<type>AE_DFF_LOW_NT</type>
<position>116.5,-60.5</position>
<input>
<ID>IN_0</ID>65 </input>
<output>
<ID>OUT_0</ID>66 </output>
<input>
<ID>clock</ID>61 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>98</ID>
<type>DA_FROM</type>
<position>73.5,-69</position>
<input>
<ID>IN_0</ID>61 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DM3</lparam></gate>
<gate>
<ID>99</ID>
<type>DA_FROM</type>
<position>74.5,-75</position>
<input>
<ID>IN_0</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In3</lparam></gate>
<gate>
<ID>100</ID>
<type>DA_FROM</type>
<position>74.5,-78</position>
<input>
<ID>IN_0</ID>63 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In2</lparam></gate>
<gate>
<ID>101</ID>
<type>DA_FROM</type>
<position>74.5,-81</position>
<input>
<ID>IN_0</ID>64 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In1</lparam></gate>
<gate>
<ID>102</ID>
<type>DA_FROM</type>
<position>74.5,-84</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In0</lparam></gate>
<gate>
<ID>103</ID>
<type>DE_TO</type>
<position>123.5,-45</position>
<input>
<ID>IN_0</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MD3</lparam></gate>
<gate>
<ID>104</ID>
<type>DE_TO</type>
<position>123.5,-48</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MD2</lparam></gate>
<gate>
<ID>105</ID>
<type>DE_TO</type>
<position>123.5,-51</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MD1</lparam></gate>
<gate>
<ID>106</ID>
<type>DE_TO</type>
<position>123.5,-54.5</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MD0</lparam></gate>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2,-31.5,40,-31.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>10.5 9</intersection>
<intersection>21 8</intersection>
<intersection>31 7</intersection>
<intersection>40 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>40,-31.5,40,-24</points>
<connection>
<GID>53</GID>
<name>clock</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>31,-31.5,31,-24</points>
<connection>
<GID>52</GID>
<name>clock</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>21,-31.5,21,-24</points>
<connection>
<GID>51</GID>
<name>clock</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>10.5,-31.5,10.5,-24</points>
<connection>
<GID>50</GID>
<name>clock</name></connection>
<intersection>-31.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-37.5,6.5,-21</points>
<intersection>-37.5 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-21,10.5,-21</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3,-37.5,6.5,-37.5</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-40.5,21,-40.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>21 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>21,-40.5,21,-21</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>-40.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-43.5,31,-43.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>31 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-43.5,31,-21</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-43.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-46.5,40,-46.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>40 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>40,-46.5,40,-21</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>-46.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-21,47,-17</points>
<intersection>-21 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-17,48,-17</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-21,47,-21</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-21,38.5,-13.5</points>
<intersection>-21 2</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-13.5,48,-13.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,-21,38.5,-21</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-21,28.5,-10.5</points>
<intersection>-21 1</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-21,28.5,-21</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-10.5,48,-10.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-21,17,-7.5</points>
<intersection>-21 1</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-21,17,-21</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>17 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-7.5,48,-7.5</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>17 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-2.5,-78,35.5,-78</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>6 9</intersection>
<intersection>16.5 8</intersection>
<intersection>26.5 7</intersection>
<intersection>35.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>35.5,-78,35.5,-70.5</points>
<connection>
<GID>71</GID>
<name>clock</name></connection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>26.5,-78,26.5,-70.5</points>
<connection>
<GID>70</GID>
<name>clock</name></connection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>16.5,-78,16.5,-70.5</points>
<connection>
<GID>69</GID>
<name>clock</name></connection>
<intersection>-78 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>6,-78,6,-70.5</points>
<connection>
<GID>68</GID>
<name>clock</name></connection>
<intersection>-78 1</intersection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-84,2,-67.5</points>
<intersection>-84 2</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-67.5,6,-67.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,-84,2,-84</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-87,16.5,-87</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>16.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16.5,-87,16.5,-67.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>-87 1</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-90,26.5,-90</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>26.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>26.5,-90,26.5,-67.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>-90 1</intersection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-93,35.5,-93</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>35.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>35.5,-93,35.5,-67.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>-93 1</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-67.5,42.5,-63.5</points>
<intersection>-67.5 2</intersection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-63.5,43.5,-63.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-67.5,42.5,-67.5</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-67.5,34,-60</points>
<intersection>-67.5 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-60,43.5,-60</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>32.5,-67.5,34,-67.5</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-67.5,24,-57</points>
<intersection>-67.5 1</intersection>
<intersection>-57 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-67.5,24,-67.5</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-57,43.5,-57</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-67.5,12.5,-54</points>
<intersection>-67.5 1</intersection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-67.5,12.5,-67.5</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-54,43.5,-54</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2.5,-123,40.5,-123</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>11 9</intersection>
<intersection>21.5 8</intersection>
<intersection>31.5 7</intersection>
<intersection>40.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>40.5,-123,40.5,-115.5</points>
<connection>
<GID>84</GID>
<name>clock</name></connection>
<intersection>-123 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>31.5,-123,31.5,-115.5</points>
<connection>
<GID>83</GID>
<name>clock</name></connection>
<intersection>-123 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>21.5,-123,21.5,-115.5</points>
<connection>
<GID>82</GID>
<name>clock</name></connection>
<intersection>-123 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>11,-123,11,-115.5</points>
<connection>
<GID>81</GID>
<name>clock</name></connection>
<intersection>-123 1</intersection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-129,7,-112.5</points>
<intersection>-129 2</intersection>
<intersection>-112.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7,-112.5,11,-112.5</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-129,7,-129</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-132,21.5,-132</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>21.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>21.5,-132,21.5,-112.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>-132 1</intersection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-135,31.5,-135</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>31.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31.5,-135,31.5,-112.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>-135 1</intersection></vsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-138,40.5,-138</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>40.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>40.5,-138,40.5,-112.5</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>-138 1</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-112.5,47.5,-108.5</points>
<intersection>-112.5 2</intersection>
<intersection>-108.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-108.5,48.5,-108.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-112.5,47.5,-112.5</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-112.5,39,-105</points>
<intersection>-112.5 2</intersection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-105,48.5,-105</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-112.5,39,-112.5</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-112.5,29,-102</points>
<intersection>-112.5 1</intersection>
<intersection>-102 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-112.5,29,-112.5</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-102,48.5,-102</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-112.5,17.5,-99</points>
<intersection>-112.5 1</intersection>
<intersection>-99 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-112.5,17.5,-112.5</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-99,48.5,-99</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75.5,-69,113.5,-69</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>84 9</intersection>
<intersection>94.5 8</intersection>
<intersection>104.5 7</intersection>
<intersection>113.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>113.5,-69,113.5,-61.5</points>
<connection>
<GID>97</GID>
<name>clock</name></connection>
<intersection>-69 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>104.5,-69,104.5,-61.5</points>
<connection>
<GID>96</GID>
<name>clock</name></connection>
<intersection>-69 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>94.5,-69,94.5,-61.5</points>
<connection>
<GID>95</GID>
<name>clock</name></connection>
<intersection>-69 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>84,-69,84,-61.5</points>
<connection>
<GID>94</GID>
<name>clock</name></connection>
<intersection>-69 1</intersection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-75,80,-58.5</points>
<intersection>-75 2</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-58.5,84,-58.5</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76.5,-75,80,-75</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76.5,-78,94.5,-78</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>94.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>94.5,-78,94.5,-58.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>-78 1</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76.5,-81,104.5,-81</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>104.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>104.5,-81,104.5,-58.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>-81 1</intersection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76.5,-84,113.5,-84</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>113.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>113.5,-84,113.5,-58.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>-84 1</intersection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120.5,-58.5,120.5,-54.5</points>
<intersection>-58.5 2</intersection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120.5,-54.5,121.5,-54.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>120.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>119.5,-58.5,120.5,-58.5</points>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>120.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-58.5,112,-51</points>
<intersection>-58.5 2</intersection>
<intersection>-51 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-51,121.5,-51</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110.5,-58.5,112,-58.5</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-58.5,102,-48</points>
<intersection>-58.5 1</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-58.5,102,-58.5</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<intersection>102 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102,-48,121.5,-48</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-58.5,90.5,-45</points>
<intersection>-58.5 1</intersection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,-58.5,90.5,-58.5</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-45,121.5,-45</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>90.5 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-63.3316,31.1778,139.893,-74.7778</PageViewport>
<gate>
<ID>108</ID>
<type>DA_FROM</type>
<position>7.5,-17.5</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Grava</lparam></gate>
<gate>
<ID>110</ID>
<type>DE_TO</type>
<position>15.5,-17.5</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DMI</lparam></gate>
<gate>
<ID>112</ID>
<type>DA_FROM</type>
<position>5,-25.5</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID G1</lparam></gate>
<gate>
<ID>114</ID>
<type>DE_TO</type>
<position>15.5,-25.5</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DME1</lparam></gate>
<gate>
<ID>115</ID>
<type>DA_FROM</type>
<position>5,-29.5</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID G0</lparam></gate>
<gate>
<ID>117</ID>
<type>DE_TO</type>
<position>16,-29.5</position>
<input>
<ID>IN_0</ID>72 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DME0</lparam></gate>
<gate>
<ID>119</ID>
<type>DA_FROM</type>
<position>4,-38</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E3</lparam></gate>
<gate>
<ID>120</ID>
<type>DA_FROM</type>
<position>4,-40.5</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E2</lparam></gate>
<gate>
<ID>121</ID>
<type>DA_FROM</type>
<position>4,-43</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E1</lparam></gate>
<gate>
<ID>122</ID>
<type>DA_FROM</type>
<position>4,-45.5</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E0</lparam></gate>
<gate>
<ID>124</ID>
<type>DE_TO</type>
<position>13,-38</position>
<input>
<ID>IN_0</ID>73 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In3</lparam></gate>
<gate>
<ID>125</ID>
<type>DE_TO</type>
<position>13,-40.5</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In2</lparam></gate>
<gate>
<ID>126</ID>
<type>DE_TO</type>
<position>13,-43</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In1</lparam></gate>
<gate>
<ID>127</ID>
<type>DE_TO</type>
<position>13,-45.5</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID In0</lparam></gate>
<gate>
<ID>129</ID>
<type>DA_FROM</type>
<position>33,-17.5</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L1</lparam></gate>
<gate>
<ID>131</ID>
<type>DE_TO</type>
<position>42,-17.5</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ME1</lparam></gate>
<gate>
<ID>133</ID>
<type>DA_FROM</type>
<position>33,-20.5</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L0</lparam></gate>
<gate>
<ID>134</ID>
<type>DE_TO</type>
<position>42.5,-20.5</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ME0</lparam></gate>
<gate>
<ID>136</ID>
<type>DA_FROM</type>
<position>31.5,-35</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M3</lparam></gate>
<gate>
<ID>137</ID>
<type>DA_FROM</type>
<position>31.5,-38</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M2</lparam></gate>
<gate>
<ID>138</ID>
<type>DA_FROM</type>
<position>31.5,-41</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M1</lparam></gate>
<gate>
<ID>139</ID>
<type>DA_FROM</type>
<position>31.5,-44</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID M0</lparam></gate>
<gate>
<ID>141</ID>
<type>DE_TO</type>
<position>39.5,-35</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S3</lparam></gate>
<gate>
<ID>142</ID>
<type>DE_TO</type>
<position>40,-38</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>143</ID>
<type>DE_TO</type>
<position>40,-41</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>144</ID>
<type>DE_TO</type>
<position>40,-44</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9.5,-17.5,13.5,-17.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<connection>
<GID>110</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-25.5,13.5,-25.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<connection>
<GID>112</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>7,-29.5,14,-29.5</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<connection>
<GID>117</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-38,11,-38</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<connection>
<GID>119</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-40.5,11,-40.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<connection>
<GID>125</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-43,11,-43</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<connection>
<GID>126</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-45.5,11,-45.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<connection>
<GID>127</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-17.5,40,-17.5</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<connection>
<GID>129</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-20.5,40.5,-20.5</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-35,37.5,-35</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<connection>
<GID>136</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-38,38,-38</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<connection>
<GID>137</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-41,38,-41</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-44,38,-44</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<connection>
<GID>144</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-73.3365,1.46475,129.888,-104.491</PageViewport>
<gate>
<ID>146</ID>
<type>DA_FROM</type>
<position>9.5,-14.5</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>147</ID>
<type>DA_FROM</type>
<position>9,-21</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>149</ID>
<type>DE_TO</type>
<position>31.5,-14.5</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID G1</lparam></gate>
<gate>
<ID>150</ID>
<type>DE_TO</type>
<position>31.5,-18</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L1</lparam></gate>
<gate>
<ID>151</ID>
<type>DE_TO</type>
<position>31.5,-21</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID G0</lparam></gate>
<gate>
<ID>152</ID>
<type>DE_TO</type>
<position>31.5,-24.5</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID L0</lparam></gate>
<gate>
<ID>154</ID>
<type>DA_FROM</type>
<position>22,-35.5</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Habilita Leitura</lparam></gate>
<gate>
<ID>156</ID>
<type>DA_FROM</type>
<position>21,-49.5</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S3</lparam></gate>
<gate>
<ID>157</ID>
<type>DA_FROM</type>
<position>21,-54</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S2</lparam></gate>
<gate>
<ID>158</ID>
<type>DA_FROM</type>
<position>21,-59.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S1</lparam></gate>
<gate>
<ID>159</ID>
<type>DA_FROM</type>
<position>21,-64.5</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID S0</lparam></gate>
<gate>
<ID>161</ID>
<type>BA_TRI_STATE</type>
<position>28,-49.5</position>
<input>
<ID>ENABLE_0</ID>85 </input>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>162</ID>
<type>BA_TRI_STATE</type>
<position>28,-54</position>
<input>
<ID>ENABLE_0</ID>85 </input>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>163</ID>
<type>BA_TRI_STATE</type>
<position>28,-59.5</position>
<input>
<ID>ENABLE_0</ID>85 </input>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>164</ID>
<type>BA_TRI_STATE</type>
<position>28,-64.5</position>
<input>
<ID>ENABLE_0</ID>85 </input>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>166</ID>
<type>DE_TO</type>
<position>41.5,-48</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E3</lparam></gate>
<gate>
<ID>167</ID>
<type>DE_TO</type>
<position>41.5,-51</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>168</ID>
<type>DE_TO</type>
<position>42,-53.5</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E2</lparam></gate>
<gate>
<ID>169</ID>
<type>DE_TO</type>
<position>42,-56.5</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>170</ID>
<type>DE_TO</type>
<position>42.5,-59.5</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E1</lparam></gate>
<gate>
<ID>171</ID>
<type>DE_TO</type>
<position>42.5,-62.5</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>172</ID>
<type>DE_TO</type>
<position>40.5,-67</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E0</lparam></gate>
<gate>
<ID>173</ID>
<type>DE_TO</type>
<position>40.5,-70</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>175</ID>
<type>DA_FROM</type>
<position>-0.5,-76</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ler/Escrever</lparam></gate>
<gate>
<ID>176</ID>
<type>DA_FROM</type>
<position>-0.5,-83</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Habilita</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_AND2</type>
<position>18,-77</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>180</ID>
<type>AE_SMALL_INVERTER</type>
<position>10.5,-83.5</position>
<input>
<ID>IN_0</ID>94 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_AND2</type>
<position>17,-88</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>184</ID>
<type>DE_TO</type>
<position>25.5,-77</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Grava</lparam></gate>
<gate>
<ID>185</ID>
<type>DE_TO</type>
<position>24.5,-88</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Habilita Leitura</lparam></gate>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-14.5,29.5,-14.5</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>25 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-18,25,-14.5</points>
<intersection>-18 4</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>25,-18,29.5,-18</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>25 3</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11,-21,29.5,-21</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>24.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24.5,-24.5,24.5,-21</points>
<intersection>-24.5 4</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>24.5,-24.5,29.5,-24.5</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>24.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-62.5,28,-35.5</points>
<connection>
<GID>164</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>163</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>162</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>161</GID>
<name>ENABLE_0</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-35.5,28,-35.5</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-49.5,25,-49.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<connection>
<GID>156</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-54,25,-54</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<connection>
<GID>157</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-59.5,25,-59.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<connection>
<GID>158</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23,-64.5,25,-64.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<connection>
<GID>159</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-51,35,-48</points>
<intersection>-51 4</intersection>
<intersection>-49.5 1</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-49.5,35,-49.5</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35,-48,39.5,-48</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>35,-51,39.5,-51</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-56.5,35.5,-53.5</points>
<intersection>-56.5 4</intersection>
<intersection>-54 5</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-53.5,40,-53.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>35.5,-56.5,40,-56.5</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>30.5,-54,35.5,-54</points>
<connection>
<GID>162</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-62.5,36,-59.5</points>
<intersection>-62.5 4</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-59.5,40.5,-59.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>36,-62.5,40.5,-62.5</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-70,34.5,-64.5</points>
<intersection>-70 4</intersection>
<intersection>-67 2</intersection>
<intersection>-64.5 7</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>34.5,-67,38.5,-67</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>34.5,-70,38.5,-70</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>30.5,-64.5,34.5,-64.5</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1.5,-76,15,-76</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>10.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>10.5,-81.5,10.5,-76</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>-76 1</intersection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-89,8,-78</points>
<intersection>-89 3</intersection>
<intersection>-83 2</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-78,15,-78</points>
<connection>
<GID>178</GID>
<name>IN_1</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1.5,-83,8,-83</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>8,-89,14,-89</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-87,10.5,-85.5</points>
<connection>
<GID>180</GID>
<name>OUT_0</name></connection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-87,14,-87</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>10.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,-77,23.5,-77</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<connection>
<GID>178</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,-88,22.5,-88</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<connection>
<GID>182</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>-41.887,-6.05238,110.531,-85.5191</PageViewport>
<gate>
<ID>193</ID>
<type>AA_LABEL</type>
<position>2,-37.5</position>
<gparam>LABEL_TEXT DW0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>195</ID>
<type>AA_TOGGLE</type>
<position>10.5,-22.5</position>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>196</ID>
<type>AA_TOGGLE</type>
<position>10.5,-27.5</position>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_TOGGLE</type>
<position>9.5,-32.5</position>
<output>
<ID>OUT_0</ID>101 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_TOGGLE</type>
<position>8,-38</position>
<output>
<ID>OUT_0</ID>102 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>200</ID>
<type>BA_TRI_STATE</type>
<position>25.5,-22.5</position>
<input>
<ID>ENABLE_0</ID>103 </input>
<input>
<ID>IN_0</ID>99 </input>
<output>
<ID>OUT_0</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>201</ID>
<type>BA_TRI_STATE</type>
<position>25.5,-27.5</position>
<input>
<ID>ENABLE_0</ID>103 </input>
<input>
<ID>IN_0</ID>100 </input>
<output>
<ID>OUT_0</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>202</ID>
<type>BA_TRI_STATE</type>
<position>25.5,-32.5</position>
<input>
<ID>ENABLE_0</ID>103 </input>
<input>
<ID>IN_0</ID>101 </input>
<output>
<ID>OUT_0</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>203</ID>
<type>BA_TRI_STATE</type>
<position>25.5,-38</position>
<input>
<ID>ENABLE_0</ID>103 </input>
<input>
<ID>IN_0</ID>102 </input>
<output>
<ID>OUT_0</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>205</ID>
<type>DE_TO</type>
<position>30.5,-10</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Ler/Escrever</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_TOGGLE</type>
<position>7.5,-56.5</position>
<output>
<ID>OUT_0</ID>108 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_LABEL</type>
<position>-0.5,-56</position>
<gparam>LABEL_TEXT Enable</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>DE_TO</type>
<position>15,-56.5</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Habilita</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_TOGGLE</type>
<position>6.5,-65.5</position>
<output>
<ID>OUT_0</ID>109 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_TOGGLE</type>
<position>6.5,-69</position>
<output>
<ID>OUT_0</ID>110 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>223</ID>
<type>DE_TO</type>
<position>15.5,-65.5</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>224</ID>
<type>DE_TO</type>
<position>15.5,-69</position>
<input>
<ID>IN_0</ID>110 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A0</lparam></gate>
<gate>
<ID>226</ID>
<type>AA_LABEL</type>
<position>-2,-64.5</position>
<gparam>LABEL_TEXT Add1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>227</ID>
<type>AA_LABEL</type>
<position>-2,-68.5</position>
<gparam>LABEL_TEXT Add2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>229</ID>
<type>BE_TRI_STATE_LOW</type>
<position>47,-53</position>
<input>
<ID>ENABLE_0</ID>103 </input>
<input>
<ID>IN_0</ID>104 </input>
<output>
<ID>OUT_0</ID>115 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>230</ID>
<type>BE_TRI_STATE_LOW</type>
<position>47,-61.5</position>
<input>
<ID>ENABLE_0</ID>103 </input>
<input>
<ID>IN_0</ID>113 </input>
<output>
<ID>OUT_0</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>231</ID>
<type>BE_TRI_STATE_LOW</type>
<position>47,-70</position>
<input>
<ID>ENABLE_0</ID>103 </input>
<input>
<ID>IN_0</ID>112 </input>
<output>
<ID>OUT_0</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>232</ID>
<type>BE_TRI_STATE_LOW</type>
<position>47,-78.5</position>
<input>
<ID>ENABLE_0</ID>103 </input>
<input>
<ID>IN_0</ID>111 </input>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>234</ID>
<type>DA_FROM</type>
<position>43.5,-22.5</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>235</ID>
<type>DA_FROM</type>
<position>43.5,-27.5</position>
<input>
<ID>IN_0</ID>113 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>236</ID>
<type>DA_FROM</type>
<position>43.5,-32.5</position>
<input>
<ID>IN_0</ID>112 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>237</ID>
<type>DA_FROM</type>
<position>43,-38</position>
<input>
<ID>IN_0</ID>111 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>240</ID>
<type>GA_LED</type>
<position>55.5,-53</position>
<input>
<ID>N_in0</ID>115 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>241</ID>
<type>GA_LED</type>
<position>55.5,-61.5</position>
<input>
<ID>N_in0</ID>116 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>GA_LED</type>
<position>56,-70</position>
<input>
<ID>N_in0</ID>117 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>243</ID>
<type>GA_LED</type>
<position>56,-78.5</position>
<input>
<ID>N_in0</ID>118 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>AA_LABEL</type>
<position>61,-52.5</position>
<gparam>LABEL_TEXT DR3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>246</ID>
<type>AA_LABEL</type>
<position>61,-61</position>
<gparam>LABEL_TEXT DR2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>247</ID>
<type>AA_LABEL</type>
<position>61.5,-69.5</position>
<gparam>LABEL_TEXT DR1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>248</ID>
<type>AA_LABEL</type>
<position>61,-78</position>
<gparam>LABEL_TEXT DR0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>AA_TOGGLE</type>
<position>16,-10</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_LABEL</type>
<position>9.5,-9.5</position>
<gparam>LABEL_TEXT Write</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>AA_LABEL</type>
<position>3.5,-22</position>
<gparam>LABEL_TEXT DW3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>191</ID>
<type>AA_LABEL</type>
<position>2.5,-26.5</position>
<gparam>LABEL_TEXT DW2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>192</ID>
<type>AA_LABEL</type>
<position>2.5,-32.5</position>
<gparam>LABEL_TEXT DW1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,-22.5,22.5,-22.5</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,-27.5,22.5,-27.5</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-32.5,22.5,-32.5</points>
<connection>
<GID>197</GID>
<name>OUT_0</name></connection>
<intersection>22.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>22.5,-32.5,22.5,-32.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>-32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-38,22.5,-38</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<connection>
<GID>198</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-51,25.5,-10</points>
<connection>
<GID>203</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>202</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>201</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>200</GID>
<name>ENABLE_0</name></connection>
<intersection>-51 7</intersection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-10,28.5,-10</points>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>25.5,-51,47,-51</points>
<connection>
<GID>229</GID>
<name>ENABLE_0</name></connection>
<intersection>25.5 0</intersection>
<intersection>47 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>47,-76.5,47,-51</points>
<connection>
<GID>232</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>231</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>230</GID>
<name>ENABLE_0</name></connection>
<intersection>-51 7</intersection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-22.5,41.5,-22.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<connection>
<GID>200</GID>
<name>OUT_0</name></connection>
<intersection>38.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>38.5,-53,38.5,-22.5</points>
<intersection>-53 5</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>38.5,-53,44,-53</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>38.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9.5,-56.5,13,-56.5</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<connection>
<GID>214</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-65.5,13.5,-65.5</points>
<connection>
<GID>220</GID>
<name>OUT_0</name></connection>
<connection>
<GID>223</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-69,13.5,-69</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<connection>
<GID>221</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-38,41,-38</points>
<connection>
<GID>203</GID>
<name>OUT_0</name></connection>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>28 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>28,-78.5,28,-38</points>
<intersection>-78.5 5</intersection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>28,-78.5,44,-78.5</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>28 4</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-32.5,41.5,-32.5</points>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>31.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31.5,-70,31.5,-32.5</points>
<intersection>-70 4</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>31.5,-70,44,-70</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>31.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-27.5,41.5,-27.5</points>
<connection>
<GID>201</GID>
<name>OUT_0</name></connection>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>35 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>35,-61.5,35,-27.5</points>
<intersection>-61.5 5</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>35,-61.5,44,-61.5</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>35 4</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-53,54.5,-53</points>
<connection>
<GID>240</GID>
<name>N_in0</name></connection>
<connection>
<GID>229</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-61.5,54.5,-61.5</points>
<connection>
<GID>241</GID>
<name>N_in0</name></connection>
<connection>
<GID>230</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-70,55,-70</points>
<connection>
<GID>231</GID>
<name>OUT_0</name></connection>
<connection>
<GID>242</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>49.5,-78.5,55,-78.5</points>
<connection>
<GID>243</GID>
<name>N_in0</name></connection>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>-49.2591,9.92262,103.159,-69.544</PageViewport>
<gate>
<ID>4</ID>
<type>AE_DFF_LOW</type>
<position>-11,-19.5</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>120 </output>
<input>
<ID>clock</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_DFF_LOW</type>
<position>2.5,-19.5</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>121 </output>
<input>
<ID>clock</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_DFF_LOW</type>
<position>15,-19.5</position>
<input>
<ID>IN_0</ID>105 </input>
<output>
<ID>OUT_0</ID>122 </output>
<input>
<ID>clock</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_DFF_LOW</type>
<position>28.5,-19.5</position>
<input>
<ID>IN_0</ID>106 </input>
<output>
<ID>OUT_0</ID>123 </output>
<input>
<ID>clock</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>44</ID>
<type>DA_FROM</type>
<position>-17,-17.5</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>49</ID>
<type>DA_FROM</type>
<position>-3.5,-17.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>54</ID>
<type>DA_FROM</type>
<position>9,-17.5</position>
<input>
<ID>IN_0</ID>105 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>56</ID>
<type>DA_FROM</type>
<position>22.5,-17.5</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>113</ID>
<type>DA_FROM</type>
<position>-23,-28</position>
<input>
<ID>IN_0</ID>119 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LM</lparam></gate>
<gate>
<ID>118</ID>
<type>DE_TO</type>
<position>-6,-10</position>
<input>
<ID>IN_0</ID>120 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID V1</lparam></gate>
<gate>
<ID>123</ID>
<type>DE_TO</type>
<position>7.5,-10.5</position>
<input>
<ID>IN_0</ID>121 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID V2</lparam></gate>
<gate>
<ID>128</ID>
<type>DE_TO</type>
<position>20,-11</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID V3</lparam></gate>
<gate>
<ID>130</ID>
<type>DE_TO</type>
<position>34,-11.5</position>
<input>
<ID>IN_0</ID>123 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID V4</lparam></gate>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-15,-17.5,-14,-17.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>44</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,-17.5,-0.5,-17.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11,-17.5,12,-17.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-17.5,25.5,-17.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-21,-28,25.5,-28</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>-14 9</intersection>
<intersection>-0.5 8</intersection>
<intersection>12 7</intersection>
<intersection>25.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>25.5,-28,25.5,-20.5</points>
<connection>
<GID>14</GID>
<name>clock</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>12,-28,12,-20.5</points>
<connection>
<GID>12</GID>
<name>clock</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>-0.5,-28,-0.5,-20.5</points>
<connection>
<GID>7</GID>
<name>clock</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>-14,-28,-14,-20.5</points>
<connection>
<GID>4</GID>
<name>clock</name></connection>
<intersection>-28 1</intersection></vsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-8,-17.5,-8,-10</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-8,-10,-8,-10</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>-8 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,-17.5,5.5,-10.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,-10.5,5.5,-10.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-17.5,18,-11</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-11,18,-11</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-17.5,31.5,-11.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-11.5,32,-11.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire></page 6>
<page 7>
<PageViewport>-49.2591,9.92262,103.159,-69.544</PageViewport>
<gate>
<ID>194</ID>
<type>BA_TRI_STATE</type>
<position>8,-51.5</position>
<input>
<ID>ENABLE_0</ID>128 </input>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_TOGGLE</type>
<position>-21,3</position>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>109</ID>
<type>DE_TO</type>
<position>-15.5,3</position>
<input>
<ID>IN_0</ID>114 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LM</lparam></gate>
<gate>
<ID>135</ID>
<type>DA_FROM</type>
<position>-18.5,-4.5</position>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID V1</lparam></gate>
<gate>
<ID>140</ID>
<type>DA_FROM</type>
<position>-18.5,-8</position>
<input>
<ID>IN_0</ID>126 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID V2</lparam></gate>
<gate>
<ID>145</ID>
<type>DA_FROM</type>
<position>-18.5,-11.5</position>
<input>
<ID>IN_0</ID>125 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID V3</lparam></gate>
<gate>
<ID>148</ID>
<type>DA_FROM</type>
<position>-18.5,-15</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID V4</lparam></gate>
<gate>
<ID>155</ID>
<type>GA_LED</type>
<position>2,-4.5</position>
<input>
<ID>N_in0</ID>127 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>GA_LED</type>
<position>2,-8</position>
<input>
<ID>N_in0</ID>126 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>GA_LED</type>
<position>2,-11.5</position>
<input>
<ID>N_in0</ID>125 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>GA_LED</type>
<position>2,-15</position>
<input>
<ID>N_in0</ID>124 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>179</ID>
<type>AA_TOGGLE</type>
<position>-21,0</position>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>183</ID>
<type>BA_TRI_STATE</type>
<position>8,-33</position>
<input>
<ID>ENABLE_0</ID>128 </input>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>186</ID>
<type>BA_TRI_STATE</type>
<position>8,-39.5</position>
<input>
<ID>ENABLE_0</ID>128 </input>
<input>
<ID>IN_0</ID>126 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>188</ID>
<type>BA_TRI_STATE</type>
<position>8,-45.5</position>
<input>
<ID>ENABLE_0</ID>128 </input>
<input>
<ID>IN_0</ID>125 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>114</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19,3,-17.5,3</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<connection>
<GID>109</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16.5,-15,1,-15</points>
<connection>
<GID>174</GID>
<name>N_in0</name></connection>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>-15 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-15,-51.5,-15,-15</points>
<intersection>-51.5 7</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-15,-51.5,5,-51.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>-15 6</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16.5,-11.5,1,-11.5</points>
<connection>
<GID>165</GID>
<name>N_in0</name></connection>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>-10 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-10,-45.5,-10,-11.5</points>
<intersection>-45.5 7</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-10,-45.5,5,-45.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>-10 6</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16.5,-8,1,-8</points>
<connection>
<GID>160</GID>
<name>N_in0</name></connection>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>-5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-5,-39.5,-5,-8</points>
<intersection>-39.5 4</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-5,-39.5,5,-39.5</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>-5 3</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-16.5,-4.5,1,-4.5</points>
<connection>
<GID>155</GID>
<name>N_in0</name></connection>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>0 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>0,-33,0,-4.5</points>
<intersection>-33 7</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>0,-33,5,-33</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>0 3</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-49.5,8,0</points>
<connection>
<GID>188</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>186</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>183</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>194</GID>
<name>ENABLE_0</name></connection>
<intersection>0 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-19,0,8,0</points>
<connection>
<GID>179</GID>
<name>OUT_0</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire></page 7>
<page 8>
<PageViewport>-30.2068,0,84.1068,-59.6</PageViewport></page 8>
<page 9>
<PageViewport>-30.2068,0,84.1068,-59.6</PageViewport></page 9></circuit>